module usb_wrapper(
    input  rst_n,
    input  clk,

    output[7:0] data_o,
    output rdav,
    input rden,

    input[7:0] data_i,
    output wrav,
    input wren,

    output ulpi_rst,
    input  ulpi_clk,
    input  ulpi_dir,
    input  ulpi_nxt,
    output ulpi_stp,
    inout  [7:0] ulpi_data
);
wire rx__valid;
wire rx__ready;
wire [7:0] rx__payload;

reg tx__valid;
wire tx__ready;
reg tx__first;
reg tx__last;
wire [7:0] tx__payload;

wire [7:0] ulpi_data_o;
wire ulpi_data_oe;

assign ulpi_rst  = 1'b1;
assign ulpi_data = ulpi_data_oe ? ulpi_data_o : 8'hz;

wire int_clk = ~ulpi_clk;

reg [4:0] rst_cnt;

always @(posedge int_clk or negedge rst_n)begin
    if(rst_n == 1'b0)begin
        rst_cnt <=5'd0;
    end else begin
        if (rst_cnt[4] == 1'b0) rst_cnt <= rst_cnt + 5'd1;
    end
end

usb_serial usb (
    // Reset & Clock
    .usb_rst        (~rst_cnt[4]),
    // ULPI
    .ulpi__clk      (int_clk),
    .ulpi__dir__i   (ulpi_dir),
    .ulpi__nxt      (ulpi_nxt),
    .ulpi__stp      (ulpi_stp),
    .ulpi__data__i  (ulpi_data),
    .ulpi__data__o  (ulpi_data_o),
    .ulpi__data__oe (ulpi_data_oe),
    // TX
    .tx__valid      (tx__valid),
    .tx__ready      (tx__ready),
    .tx__first      (tx__first),
    .tx__last       (tx__last),
    .tx__payload    (tx__payload),
    // RX
    .rx__valid      (rx__valid),
    .rx__ready      (rx__ready),
    .rx__payload    (rx__payload)
);

//wire[7:0] tx_fifo_out;
reg tx_fifo_rd;
wire tx_fifo_almost_empty;
wire tx_fifo_empty;
wire tx_fifo_almost_full;
reg tx_full_ct;
always@(posedge clk)tx_full_ct <= tx_fifo_almost_full;

usb_fifo tx_fifo(
    .Data(data_i), //input [7:0] Data
    .WrClk(clk), //input WrClk
    .RdClk(int_clk), //input RdClk
    .WrEn(wren&&(tx_full_ct == 1'b0 || tx_fifo_almost_full == 1'b0)), //input WrEn
    .RdEn(tx_fifo_rd), //input RdEn
	.Almost_Empty(tx_fifo_almost_empty), //output Almost_Empty
	.Almost_Full(tx_fifo_almost_full), //output Almost_Full
    .Q(tx__payload), //output [7:0] Q
    .Empty(tx_fifo_empty) //output Empty
);

//state machine
reg [1:0] state;

always@(posedge int_clk or negedge rst_n)begin
    if(rst_n == 1'b0)begin
        state <= 2'd0;

        tx__first <= 1'b0;
        tx__last <= 1'b0;
        tx__valid <= 1'b0;
        tx_fifo_rd <= 1'b0;
    end else begin
        tx__first <= 1'b0;
        tx__last <= 1'b0;
        tx__valid <= 1'b0;
        tx_fifo_rd <= 1'b0;

        case(state)
            2'd0:begin
                if(tx_fifo_empty==1'b0 && tx__ready)begin
                    state <= 2'd1;
                    tx__first <= 1'b1;
                    tx__valid <= 1'b1;
                    //tx__payload <= tx_fifo_out;
                    tx_fifo_rd <= 1'b1;

                    if(tx_fifo_almost_empty)begin
                        tx__last <= 1'b1;
                        state <= 2'd2;
                    end
                end
            end
            2'd1:begin
                tx__valid <= 1'b1;
                tx_fifo_rd <= tx__ready;
                //tx__payload <= tx_fifo_out;
                if(tx_fifo_almost_empty && tx__ready)begin
                    state <= 2'd2;
                    tx__last <= 1'b1;
                end
            end
            2'd2:begin
                state <= 2'd0;
            end
            default: state <= 2'd0;
        endcase
    end
end

assign wrav = ~tx_fifo_almost_full;

wire rx_fifo_empty;
wire rx_fifo_almost_full;
reg rx_full_ct;
always@(posedge int_clk)rx_full_ct <= rx_fifo_almost_full;

usb_fifo rx_fifo(
    .Data(rx__payload), //input [7:0] Data
    .WrClk(int_clk), //input WrClk
    .RdClk(clk), //input RdClk
    .WrEn(rx__valid&&(rx_fifo_almost_full ==1'b0)), //input WrEn
    .RdEn(rden), //input RdEn
	.Almost_Full(rx_fifo_almost_full), //output Almost_Full
    .Q(data_o), //output [7:0] Q
    .Empty(rx_fifo_empty) //output Empty
);

assign rdav = ~rx_fifo_empty;
assign rx__ready = ~rx_fifo_almost_full;

endmodule

`pragma protect begin_protected
`pragma protect version="2.1"
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="GOWIN"
`pragma protect encrypt_agent_info="GOWIN Encrypt Version 2.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GOWIN",key_keyname="GWK2021-10",key_method="rsa"
`pragma protect key_block
CjNoDkJCN4W/BnJoiMP6blGJPezm+PpHAZXzHOz/tHCFN6ukE3pn+Af5nblDjtNDoFkI7XIIny9l
rZLlkyR1iysgazFvL90JUSImK867DQ741LUWFdB03mivQ6AuoYJ27+v1lAF9sSSBSns6I0cErz9F
cD+Le53jH9G5p+yTwE57/EXRHhH3rhuP0/HqwbOR+OuWATAuYgLa0NeG/g9pz0IdjsPMlzmA/Zrj
EOcVGx2wDq+tmDYadtb5ru6+luW2nsH+WfL0DGvWP6pnnpf9nShtDTutFSp06hiVxZXJSfB6hnCs
SgCir3R/9CotfqWHcovvn9YJpp3AQUi4HaaNIQ==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=31712)
`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
yJgwgquD9t3YhJk7JapAPPdeshX0dP5+l2QcDwj7XFLVrU3ZYymWudbSBMDlBTG56jJKn3C2fARJ
8H50VdWMHC+PTG3C0ye2FOMRbNiOvz8tVqt3cBP7iVKZAmYgaLVwzyXFr2zV7B83HAEGR0YiD9U5
VKbLLocz4NQ2VZFNGjO+3ofZ22ZaFQWRuwbBzKxibDURhNuFGB9qZYKp8xkcbkF3qbBzV795/b48
ED92OD+FeY7ZhtIcdlzbY00ATM6YRhmh63xNkrAZfZzwRpkxSMKkTVEcGK8kPCmBzGO65P35gVSb
YhAERYeektBOZkxcAxkUZE39QocYGMxIplrVy+PEDmqENQgH7jCiglhHBPlu6V3Dyd43XEZnBtEL
3lDXp5+qY12xZAll45tWnDl4kZVbbWhj0gSUq4+ZQ9xOygp+BF+CITX2qYDJMz21/M3EVjZNna6V
tGtdEATRmNhoFszbaDHX3KdJVooztNUpYzb0sHjBLqDVZvziqB8KDSk3aTavHZUT5hcGuJTOTFh5
uv1NtDMm5NottcU79uSB5d/YoOL4TANCQRipd4ZBhCapJrVnjNkyqMCA1w+SBSP5M1pBJs+tfKnQ
KTfbGGeET03mBXHAZv6xbp59Dw6jkvIZX9431KAzMl2Z1kevNRO947bTLcmHWx5BElPxoJli1AAj
pZh0EDNulMDMyZw8zhMbg2L55t2hdHWOZUOBYDZo3a4vPmfkA+XQ8IeEDDkpKxopL4c+KpX3AEEK
aqH3rc6CVARyslbRhN7wlK0VLeDNrFkCUvhwX0WSnZUP4VmSMccxr56ExtadGz8/P5pXxAmbUcWr
6jU20eVkbPS3pggwal1PrtmxNnNHbrRWWN2M056madeb78iuW75uLi2/vAxJlcuR2fEQq+znKoMl
K05ThDRaMYi2x1aWEKs0KCnGfXqMYoy4TTiVHESrN8bC1tSIQwm4uJ0WFBWsjwr+gaslXMXGgmj2
aBhBu/tyLvzP0kjlpzDvnudlOiE+5j61M7y85hmhHXIbUMueeLenrgJ300QMruX6RSwsGzFvVfU2
SrBEsMYRDlxIpHizYs4LBe9x9TonlYL0QdpvdTVLBsbgc947pI2czKse/2eDp7RP1Nls8M9T1g9a
kGiis0kB7IRPNtVP+uLEBDdo+4nkCxyjASHjZzpqhlji8op67BHcCUqD5ZE8FjRylEQz/BNr5ryJ
yVwtysZygpWwcmMo61Jix8ZMvYvksgd5V7iTd55x9ZIZ8iH8GgMA9YOGAu8AnCmBuePmm/MIi2fd
oZ5UcHogyI3ht0+BUJIumDirYwOefE1uVYC0umW9wOqYgDxG8sN6whyUL87IbS4UlU1al2haedht
sbfUvwltVAPkx1BqqswbCEvtYLyXh3mJ9Uiw36WZHt1qmg/3l623J7DipNTCI3u0IaIvVYPhOcuH
BTB819NNDnczwtGxW+nrRwB9E/5qJOjdPSbU4kPKQR8BsHONORksGi2NYaROAJgEThMOxy6nPv1g
VtZfviAswyDgBCoQc3slP3RzN2uKgu4czeiyEm7SXhkDfG5zPM4FFSCdGWiNzfIq0hX8d2K8e4If
LB6vNu5nSQZKPcKuPYXDDqRuRlxsxVFdEG4xC92wdR7VFEtMH3TklEiXidmYCLpHHY2Xu0EFrW+1
nr13U8mwiVwBE07uuzbZdF36tbx1rozNdx9w5CT2+tv5P3LgMWYaVcE9I5wHmr8nzsaVtEH8Fs+7
PY3M/6neos/A6ot+5LhLsTspC0ndZn3RIZKWOWfJyEYWNXrR2YnIvmrJ7PE4fktI4WKWbXxRNgpW
rpPHC7sGYi0PlamKlZp20TVh7xSkOzc3fzBgW6zttG/F6VZ4THlHO1YYcPeJCLST4/coiT32MuOB
HEZNyK2Jc0p43pGpEAu3dOJmO32i6naxgTWYWpwtDTt2ygj4VRbRyZJi9Bka0b8vFmHETRF1sqDj
N9lvxQDYXIBfdJIClsarEZ00xLWos2UNeV6HpLGsfKKFSaPKjwrmrXvWmu4i9Azyap85eDa9866u
KnJA7pNwE67VPH+6i1uEqb/zXz3Xcol65A1+6pCiT3Yu8eBo8RKi0KikPEw+66noZrelJqtpu2u5
MWbHNXY0hdOSMb0U3rl2WxKVCPLULST+bNT2OIXxQ+Xa0uorK5L+aErWxOmGYssakYIhI02Dw5/R
DUSlyYs+5doj5qMEtmf0TPkddGiYjkLtnUrM/lWIbcY/aD2giaJNOKiExTuB5711kar+mNuZ44SK
D/2Y+Q/rei+mN6N4BPgUh5Iqhae3ewxiP3GVdHHB5+UZiyep/H64GtLHeRWGv+Xuf6YIUeYMH7Kl
C1fcBYwKA96wH92qg07S2A2fe1NMMu/64ipW/1L2+llr8a2JfPIwdzG6U8jwtAHvISHHIe+uKnxk
rQFlHt5uTnvS1f7mvwrZ10dUe5EMm+y41dxJW1pWGRRAC46ToC3+C+3kRJv2TyURu/uAphgPr+jz
QqJKMuxocLk87b7WPnCcbTD9riHNmfPUCbWvMqEZn0+f/oZOuVHE9L3JX5WANuCuUDAXBgZqf4zj
Pe152OG2aen+e50dPWsi+X7r1oNkMf3Rh4hO7R2yQmJGy+FGht7KeYxxBFgsPmJ+8h7+0BIO7rep
fFsS93wafcYqCXMJN5OdgLr2U1jvlAYHBtpC65wHlcQyxMPNdKfzMcZu/IFsHF5NzZcLGLZXrKFy
OcQiratTY7KupYByF04NnItvVfgMAg7cffQRlQdot0v78zDZ03mfvM3YdndEFtpXT0/fJFwKvm16
mqVtzYC/3qIhqPSUpl/PD7XXKOsGWFuFueTFtqc5etneGZe7x6nfLN6ebIKDrw1FqVQ14rZEqLux
aBheVeAVoW2DvVfVq9camVabOjbFNaYmB0jA+cT/8OFpXledZ+HTsrTMVkeTQ9llder95W2wFiL1
3MOGjM3rw/wzaOTWg1W9G/8wkbq2nw3nCAvgBfoWciMzENn21FhOkQA6EpoBeMbnspJjKJ7V6JsZ
ToLWYAfgtMP8oO5uMLiutUtkRD9gAftHiCW+9xjQV/FJrONM/48rg8t6Hmv7f7B1fKrpDXcb0V+m
TyDAgolDb4lAba+v9y4FhnboMVmx+gBigdbrMTrRmgjLYKiz0Lk2o2ZtGWlXfRJrIN2VIeBQASwt
yFRQZ0VGreu6cc3GbIK3LGi2kFbkrOephlNs10IdxBo7TLcTpZMTDa7GHLbJs5nTDxJ5Ou2aIhgl
grvGzGS/8l9YtsnfAlspbe1qEyhPQl71x30sS/mQ4bSs47ycCQDupJ2hmR3I1zFl//qW6/sgVKNw
bgZgxEQqqTWQUZFAMj4FeIijYChV657ANfbNw17ItqMwtIVzcAzWvouA28o+Snyi107XYqPnLZ+A
62zwcnA3bma/7Sv+iLqPAwVyUkeA/CdNUsfvycyGVlRPvQOijOuwaHBQ2mpNFGiyi3izc3IeWhQx
WpFENZiwtMxOQQ5/DR1WdKWz59kICr8gFC2zpiphsZxNf52no6AyGRdwiPQKpyXVEDsbkiq4vmSx
oyBnwAwUOy893i3XJZ3J5++MapPoZlb4C4l/DyuegOJOZpR4puMa76sZZXDePfkn2g8OM17xxLlB
KTQEBDivTZiT3zzH5kxJGFVXlRecTRQv2e337ihpAg6COiggi35mGWaSDbpxJt2w0Vv6pOEbmUDz
sHx/9/oWXS8Ci5UblooZYN2hN98hL/dxfHpQ3S+9WD+KiTAJ2k5Xu068fpb670KKGHpwd1Y7R1iN
qO/Ltzgv8+Fqg753LyQP1ZtaPy072onZ1u0xgtUCIHKugV8Ojcit9Wjdkz0JTHj47mr49y5sB74R
byIlTHt/bEh3KxcXnI/24lTPmorKAVgYgt2zwMnTWLBjYH+yL/Uq50h2edfZPO54jp9+3MdGqLFl
9KjWc9SLv4ZQXTOKzydike8083wweSRNZCX6sDLIXWkD70EBrv6odu2kdnRaDp94NMowGXdrqtgP
n3oXIuMwnv4K9dvWlbPZjCyeTn2qi934MLeQMTRkvT1K6nZ0Hf3ChmB4nFc/eC68ACF7L8PUb/w0
GrxmAH6av5z31GkJ5FP+1Gp95u73QwynzW3C4dgFu/7njmD0byLcFwqo1jEMxK+O0lXq3hFKw+q1
FGsBPKqmIM3x/WS6H/jNqekHXoxWr1Hc1esIc8eYBChccKxsTj3CxN83s3FL80/XBmZeRcBSSJ0y
JSoIXddc9I1sxb0Pp1Np1S0jWp1Fo8PRFBf1gSkAZLWzxBLiaobPZoyZj+TqjfQCfBKCX3Fh5qGW
dfRwo4AuiLlhEvzNY9VXaii4wZ4CySCTAl07LcykfZIl2vvS8T0LKsPWiDKdjY4Qmm6N3tkr4acZ
6KCU6nI4Xcv5wIf+PTLMQIz43yR1O/RIuL5cWuYiNcjNMV/RM2kLRx9DAjZt/+53uEIAtyHCdFER
MDF5aDDOeMHBEBxYlTGtgqPQQSqEf3VUvfHyvfB+wp5GG7PeZGTBPc4D50rWdbE2YZrje+aZ3YjA
+XaKTnXEODoRlSNpvylkiJkvPb0zjEX9Z0vSCqZtoeSIkZepsiMYziyDkmelD5FkQIMmEZp3+t7c
0O5DX/zPPWmsSHLNOBALrtCfiWTrAsELAoYIpv88T8hmeYxGcIcOczSrmmqlgEFTHrbleHZr9sJn
GDKzPW9luGy4j622+JytHwvtN0xm2qhMFdBaZH7vDGVqpKzxHveFqNQzsXwFOb3ZH+FAdTD//XjI
zvN/uaYcOMp5KH07rUv8JfTUvxmMMeLN0EURl7XzHFi/hTgfoIqjQtTgbZbGxBwb10CFhFwkgaS0
6B23vhewC4W9JwLas0IfuXlIOpqbxvtu0E2PIcaUG7HZMNaB0moylxOcvADx9TFieSxCYgQXr8Gc
oI0gIUqiYMJm/wGGb/qEBKSF9sJ+z0ALcjHT4SJR23rLw2nx6jjs/swuKkTIjWE60PTn1QCVyf/r
i0ycGX/zr7iVjxJw3xTCzWDM9hBvyNgnjroRgeRgzB/trEapbJ2kiLcvf2t88F7fJG1/PMTE5xf/
UeEdAkW4eHVTtzub+M3fGY0ijfPRNFprX344fJaHh88mSOq/HMCJJHivuiZuDf4CR6ulspErokAs
YkAOpAu6t7x1sVHorLAtEWTtFCW3ejVcMSV5yzCCcQFjPXVWSfj02UxMpy7MjYQ4NBwwWJsCggrh
zrDWTGMsiyBNTz98tVF7UeQBs0elUbJpdUcp5QAfjsZiRJBN1dHsU/BISiExJv23Rmvz7Smf6hle
ygM3A5FZjvT2JG0lL2FmhhWibKROG8zRcHNAB5XxWOzb7YZ8Mf0ArM9dFtWf7u/oFrdoA97V4dY/
yLbhR2bjgpJzZCXekMxgYrXslMVteTK5/1xuMTZWuOtlxLqHgjNvJdlriH0I8xVKAb3aW4FfCDYV
ACjSaw3pP6Z1Bznu9IQQfscBFNjAfjIEmZESfu30MHZX/7LT0D3x1mMtdO6tt297B1Rwn1i7CSy+
vQ9qCYt7RoOVJLCnee8i0FOLmy/esCPgt2WB3b6HUi+Qn2OD75vkW1m9I/X2dN56sFNRIl1i576Y
zEDdSHyXMZmpDmN437s2LcCiORoALc3x/Yg9+przXcrpC3yBdfu3sNqdwmlV3FLyIYop8sEzFyZf
LR/ZbcngQgGBQcz+MM9hs1AVODwa3co19KxcOI3ctnTJZB2ZLl20APTpP1GsJnjDG8LUl4HFqJ08
QqNYLFwetYE+Y9iiwBpdlAGuqIyxDtE6ABSHyWv1plfgFHev9TonO4Gy8P2zc8io7XrX4ECTavWU
0Lb575gnO/rbKn/DY57tHr12JNSo/7LRZdfaAPNH44gZu9v8ZyaodFtJ/wrj5uKiq01vHNuLzBfH
f9DE7c5vIzHo4DSUrntGiyaiMT7kWzzRwN5BIIIRz+v/Pk/HJS1UHTqIRbluax+nckkA6v2/VJne
4gRNju4TLELy28Lp1O+3JvHD1Jfgpnky/U6/ykh8Uf5sMfAwPRmjmt2evw6igZ83vJkH8xlEfGSq
xkrrH7XvXfQwijISnICUapSY2dd1jshWFuYu1TNsOY7uja9f4SymLSaPm/7Y678ATDzxvs3nlusi
NCn3agLlnkZaYQz1lqTJqz8ucVmiD971BX81wdcLjetNmDCVJitUpV/kBoeZPOM7DfhuZTFsb+ii
7hslJq/IFsT6rNyh3sZKbRS7AcwTChkZ70BZWzzE8XWL3uy00IZAsR5HohB2rqvajbJ+EUwxrRWd
/0wDJp0rmpDMY/blTXrcdQ04NG5+Dm/+7F4rMwKDvOqi/U2df4MsggJXEoJlDeufGC0iVq6BDHJg
+8wimQHdUoPRzKL0pJrb9buY6d+2x+VySVs/g4sbnLr+B8KX8q/8GTEVsQvBrOm8US3X01N/fDwe
J51UhvOeKd11HUYO5AClPN9wMyvtZHZz8G6JlPWXjQbUUOztSzCTks/0oY0KgOpO/V0qBBrLT1Hm
KEH6q2WFbw3fq+JBwZvp22C4npoLf6BpapTGvTglWItOdRB30wCOb2f7iDws1F9KdxU+1qcyYwOP
dxy6xs0OEkxEU5aDFyNh3daLjqMUJUh3GzCA+CKRm+m1380T/CxNJxhYbOd2VOzGSCJNbqmUVAne
p3B7quGEyhaNh4/oluplQBVgLMcN4EZj2tJpJ0GYBhECsD+fm7pkdb0tkel28qgXiNFGNNqTJgiB
2jfad000iKwymCDtXc0b/JwQvqvuDw2F6wVMEQtVg7+V4UByajeyUAiNlK1QbgVZ1a+TUU/6Sq0f
MmIjFzbz93v84FfRtZ7Jz14xusOvA2VXJW5VM0OZ2xBMQVupGQQrAUuFEPGfb1ZKp2XGkJSdOILY
7n2UMnEk4iOUo60CYe7o/PzeVO3WOiXKt7k2cpcuY65i2CzUnoZuOvaUrrd8UYhCxv8l9t14+dIp
mYV8tXmcscBRVOWUebA3ByiisyYVx/EAHDyNJldJB201fC4Zp0SPylT55BOllJ3dvTR8jamQJiUJ
DMf1K3o2eNeMeS8Rx6y0dxEZFs0HltgX2uWEQByR/Fur2tlTq012GCOm40DX9MGEd+t6mYCbKEZP
YpY+i3OQg53xOUpgyahqyAn0CIuA+ykNh7FHOYmhSbcBSqIM4xmPTVGpiFp1dnhEJMSXeFoInyE9
dRM/Lw39uQWMXH5K8G+PZI7cNlm7ngS8Yo46tXOeC7tCLcLHNdt/zggpUfEt0BkynlgnsY4Bjg60
SToNBOpgX3mYPEkTvMJtoCaMu3uEENUkbSFaphI8oL9wk/f4rvbQEAV1MzhLxtj/G7o8aXtlvmVq
f4oqYSoEZb3Zj6U75ZBBEDIUXDi+O59S2Avd+hYvZGL93Xz1cswsx0uR4SFF9dYS8hwwTz+95MXl
NbilhvJsjY/cQcg24kaSA+jH1Zx6TiZZglw1eygOJk+v6q9hgUSByT8o8sZChHVHmqJzX8Uf5PSw
lsFsalJD6b8gXn7bBoPFmY15sEnOPuy5fsafJo0mQR1Fd5rtDycocT6sakE/POV1ZdsaRl7FopSZ
z3Z9QjNd8K/A5Jn6cK63jAZ6LEXLnyIZDdXrI5IHqJu6+IJGdp8uvTIs+mHlCBXBxg/V8UAINd2A
20Eb5UIx/P3QPNey6TTkUchlAQTN+syoMpELP4rIfK3fJfRlUFNFHz9qXK5tbOY9xOgzLDZZlYZz
16ZhqIwXrvu7vERpqtL09co0YXaE7WDCrN4QqteATB4rdozHtdbpaJYcdbzYBQNflMu+fjnY9eIP
C7efCNLFnf/bpkbZa/fLU8alr1u+ocuE33b4xYDSPOwR48lxt6jI2BdgBp/t21/kS5dL6lQnCACF
rNH8EF7uADG2wzbKT3AQ2Cd2xpDssunHd33TPEx9T6ttwG6HNaHdNwn0GZC7kAT5nYmaXdK6zR0+
+6RWgDhWr5bkWmqs4CVUtH5Nvk51CE4z3ldZfk2TT0R8efud5YPMqUKb1+DlClothTqtkTX8IYEF
+0FICiRlcJLeQJtCztFvXuAsc4y1u+Aj3T/zJ55V6+AmIqY4V3kvBMYLVrZPyOxH3dZKPheB5nP7
HP2ZXcH4B2f5Aj2YbMNYXyjzcQ+OC0rTVYLCvwEN/12RYn7gsVmi7gjqP9atogf4pUDu4Fp7loMp
hGjzPvZa7dr2syZECfS5k2S51cqlHD4k+OAX8MXsVQTVRB1nZBo610CvlUcCHDqkshH/214Wa+wW
SFmUt/gVSNH4Y5Xjh/Y1l/Te9rBkhucReUHrN4Ixk4aHqj6vPXd6E+K2+acjdL8jJcuPWWtDqTex
uAb9xtq39PMsday1cVE2ApXAqpNQS388A2mAtgSC5GCFeGzX3LuTYt6oC644TM/53EDI6pdrqhaB
bQcieUKD3i0hX+gbCprq8qx9d+gg4WfmHkeKAWMdOFpCeJfwMJS+46V9lwESu9oRr5HDMJ3nxdSZ
Pou+ZBArUpj9DibUo4p987NbPJL+ztMfU3cGKBsozsOhexFQti+7T70CFzLPEnLbO04Fa8BSiDkB
agwE3UG6BT7B2ojkGc1kPZPaYmzQ65WSMhBaPrAZP0jaGPJXssWkLzc+qgQLy2pHvXFgSpBVjhWE
R9YljMPHxjDn7oawrIU0PB3x0Qy6hu9iNot/aDvjs2J4+4eQDDS6F1wAG+ba4GGqsL8Cth8gBxIe
u7UxPRCXQabBxLm8/k8GHW0rGMO3S6qMfLPAmBwSXcUo+Wge4KpsYHkmr4VALwNHShYAcrexNs8F
aJt1a8DqZmXtP7xEmfU/7/u+9MkoBOB4yXK4qn/Glh5rPY8d6vWJj/rJh+2v0a2/jBtAkjKztJIw
eYIt4PrhS0lWDInQVC0PJtJvp5EP3beAoY+/Q2lTwU6pLdtPeRPRGxWdPut6AT/RE+evV3UYPXyd
dCCbkzqtSAIka7l1JHURpZ0VTb+SdcdZ1iX46A2wiRsp1TEJ8tDgyUDAxFTVYCz5q87FK9zMac5X
By6UzgXEtUMk0OPuzD45ilhQUU6nAyPYLvVQcPjMRY8CDdwyYcyol/a9/lqwGziCOFKm0mMvjrq+
Ck4h7o1N17jDPEkVWKEk53OgWydy8qy/lcFCLbjX4OhPKAuiRkO0IgCVbyJWv3ZX4Os7WTPhER/Z
ElHMmBBFmsSoTY0xi6uC4GZICSapv7LonNJycZchxd07UE7zj2+ywIoDCYU/dyT3wdVXFuy4WvvG
secrDHSLTTpGSf7AXuw1b8AEfnwX3A3jEzohVCoosL2pZ1cx8N3Y4md6yNFw4AbTpKFIdiDb8gL3
9x+VritIAohjpR7BQfVLk9jRcNRO6y0uG2blcNyaCcDmrAHEoqHy9O3PLkNttArR6qG4OWAr4eIz
4tG1Ju2pSE9xlC6sOeV32SKytFgIACwfzyYYZWmCoXzpI+9J2/vFXIQSW91goakLmvsIYIcElvbO
JC+sOsjAiLWNXqvh9fpBXoAZauOXWytTo+lRcVJF3YQY9cGUsO6zcUEy6J3+iuyeJHebae+ArFS4
fkfxkuEzZsMFXKFLJKOca8Yz5nOAh9g3hX6U2aq9zwtXd13cCTdpkyl/6n1eZjQFQlZ4AT+1Nek8
WiXj+VCKZkEpmofyVYzAPaUT3MILuyF1wPuOPt3rP8PzcyHmbebH25piZ+Q4lPXcAILb801t8C23
SZBnfbo+vKYQdxBb5YcQ27IXvSk6TJ9dxha8T2XoegW6YZJX9K1KuNmjMEAyCSda+mfRWisJOgjr
SGIXgGFggtoAZDi336oDdnwFdD3tC4RWMRFQatDgm1+ov9SwPSiB9EWLyFt8alCVgBQJqnJf09pj
xsFrA2VuF1xaLAqyHEfq/TLE5fJ8GvcFhIMuZLmVahIWvbbdJnIAaDWFydNZejQ5Z5ihHNvXJNyC
q/dNAWL3mfbV/uLz27xUyYpLTNVvwycUBDImSqosiCvWQXDkEQE/RhZqL/1nLbpyigSWPleXMSae
fVgvkjKks6ljAirZtuIktb9kwAigB8+cjhdYqZy9AogvjmfcpCL0iO4yfyxGMsILUienjsER/gO4
N9SDKvSJ5Orf/GGI6A6gwepcUPd0a7nPtGXBNiUDElOuPlMfN2uwoMbvdfm3elQKau3lE3mSUXgI
D115XRyB3n++W88TtIFJ3IkJazl/O3YtZFbfjmatb8vD6ANE6VcyPJtA+ZZ4et9LtxLLRA1Cn/6o
pNUbpzPxfciP2NmKHIOC8jhPaoIVDtRBCpW0SbhYsrCIB4Xaqh+Db7n984bzJCmsL27113hy2cpV
93mld3BI06gomxwdxW6DVTbMrEJ7dUKWpEIfnLZLtmYvqnDktkUdybcFrj3OCKqzlOb/4pF6JDNV
eFStm9bRb+0V9taSCqpg0owATiaUYywXuGivyVg9IoqoInnji1GYhbp0/UdH0IiLG2iyR7hsmijT
1BIK2PHm7JpzNibfzzV5jjmWE7PUGOl61T1oyMf+R50VYdCIQ3jZVBePTDbNluYb6TVbqZyz+zdI
8XhqWx5COJwsLBvP6wRb4gClyPlJ/pJsVH0lGmC8qXGboWyZeYyMf7A1TwsHhBnbMZehl22tiSsf
ujOwAP8jWeuuJyH3z7S12OLNvGuex/36c1Haom429JA0fMDIa4ByVGGvauKaA8ALGm/qSbHiU/is
BS5SGWg9DRe5NHPFakGt2rQHpIwMWOubf6XyZzDDt83/0QX4tyOXXsNKb0Ac5ib8M/bsCX17/ti6
HlqZenfgjgQ5Wiiosiw9vOA6HpicZA0g2oeTDVjgSyY2+m0rlXJFSm+RPw7dwVErH4drDOY0BOdm
yDF+A4ewut/ij1veTmYYysMpImAcZ0JBcwyntJnDkAWBmLojqyLoE3QVxBHz0zmKnFHdaNoMUXCa
//Z4dDWnK4rtKi19QeqoDeCHl+TfY7U+LharXsLWnXcnpRVFA/XJW6qtKLVvKiZxCJHf7t2eK9DG
UMzPCG/+Npg0s/11I1ZPaBNclICBzTntM1R4jggt0n7nlxCqtVlfCvovs8Bbee3ew08sdYlH9Srm
IO1j0JE+vQRX6EMZywi6/uRgUaSp6b/priW09LdvTDq5gvu+VwfBkbSxt9zZVARjaF57bnu2BRzo
gP+NDkh9EG+X7vqwtMd/7bYizFy5AGULAilhxSidutK8V0Jm8KuSI3fUqdC86CJaO8fcSdwdVLxm
lEBpGcl4kYMumqXDD8yWAvGBiHd9zbdIBzRohSOP8J+8H70paTS/AEOXXMDBqlr7YrypCYALnz14
QAh9jLJDFGvgA1QtlyHzOflLAjKDwyCoBpuQS/f0GaFWoOu4jUk9AApkyTvEOOVTElOWJaOgXRDz
xTdjNXSms5sldyBFh7SDoIzSpZXaZ7qry1A/VGTVL2gwZc8tO8hdmz1Czbf3ssi80JmTdtcCTeBn
NIPQmYcatCHzAv0a11as7i58af0dXg1vnZFGOHUj9iBVHWmf6V0veoGyxeTDDYP0R906eDA3eNE1
499F5QFglZ3ziHV+TUue9c008PDw9LyAE7DHZBowuSbafH8FZWlYY4tOWn/tGQoFalEeEbs69wF/
Rgez+EEt9MDbN4WaI86E2mlM9mdvWgBRa14HvH9ZAp6GCSMcMwFpl81KnghYEySQY9GQVKb+CCdN
cioSIQiP++MZ7GowYRA2/oRY8BPJwRThT5oQaXPNhQ5UycGH0ZMLXKlgCflBpsUqnltPEkwQxyCS
m94k4TN43KaPx++9iPu6MjYStip65jcULlM8xWO9TI87o0bAyzUOaFfvYISxgJN/jzklofVZDuCG
tqqWh8aDWsWUwkEmz6N7zjVjiaWfpWO8gDEqrquNd0TzJJ83wD4KqrxLkbW3XP7nm0ks+tHXTeb/
iuUR8PbSKbLzMs3PSXK0fz3KNJ+4jMlK/7FnCCBHErdvfFcHwyF8/f21HfWXZ2Qzw+ehmKgF+Ea1
TTQJpy8MZc9yqByLKdDZ0s99tmIANj0bqWjmEuDNtoAjO44CSn2/F2RaZnZ5/1sqIrID550Ucl3z
qiKOzPX2rnAvujFtGZ0Y5z6Zf398dU881fS4Si5mFugNEE1+Jf7QwYP3/UYmPcUWsxj0D9YummKC
/rouOU0a3b0O09hRynSvAyg9cV5VMJxcxvPlkWcz7rz5/TVLnIw3gK+9+WGG4eA3QKry6uwRMIRk
Y3LtC6f3Sd/OIut293I9F+jbl9ZvuiQxtcc+cbE8x+7wEtyMEUXcFZzlbIzAFCsnYV+coLsrSbiR
qQ9dPY4yUZNP3Rws5VLJXe/2ZEFNSU/DZd7sROPVtuo3I5MxmO/oXJmVrwXMmiqbv3tV8zpfmmBQ
1LEhmRYxZt0fxeWFWa5KdJY677AA9XfUJLKXQ3NQpNUOJgZ5m7E33RdS4JsipZm+6nayz5fXBRn4
TXwNnvsLMJAhILNSt+lLtkzgTi4qn1JDCVuLns+j9bIbjKBiMh1PHTN8rtGTGpZuw1jDt14KUTHN
3AsIIM0NGbWaFiWWfQWHeJ6qxNQiHMS8zl2Tle6Ee678K4WWdz7D22ERKDnFejrLyAivpp+V6CYF
BBDZol/IAVcRhSiyuG2dsKmA/QFMwKnW801DMuxDorYnvHHofy3bxGVGkBJ5S00F4bE4D8zKM0fT
g00epO4WTXuD+UjRpp7ucLaMwGTCxADquy1OUuJJ0XsKxdI+aGze9godqE9fw6BsmVx08SL/ApOK
znYe8dx0Q7xU5Zo0RV6zhdR5M8sZH7PZm5QC3DgY4xKE2lTDuMxghKDKTSl4aJZz0K2kJqqjpun4
y+iPv9GBNKV2yUhdCHvlg6WJd6jTNoDp2Hu+UKByav1lr8PMTYP3IuBYPie0pBBAgMuThGPG6oTU
XOB8cQRSgunAB7qrbdS6dyzVUjpO4UzIgXjze9A3ww5vfjE6IlBPuUmlmNzm0vNhFzdF/xKN800d
Nt3VxCHmfmOx3N2BuhKqLEMLy/wGFmFTGxIT0Pzo155DB7TBH3cxetXDQMecS4BRnw3h1Oi0C0Zn
wRgmfddcxCVz2RNPlt6U1CQ7uKouvp2lXWakumeNGvCnMoQfP8IOqN6kRqOO2kHzTG8WUilbQD00
/Auv9+348KOPJs8gpmqAmHCzYvsyU8jqpa6v2RuPAoEGOT4TqsXQfLHon1idwS9DarDdjQLpdIBz
ICZusZ9102W654mI/8Mmwecm72y9Hm/7+qOcJDko4IWXXiGmtqcM/BwQJoj6NQf/8kcPmJ7xSnGy
ZFOK4lJnKKRxzqQGgYmZ2Ff0XDvmD8cHzgePsTi6XbWt3+wqGQzHx6gw1UdmACBJmWxs/GEZr1OS
Z8hbc+B5PEo5K/I1JTkUPYm+0vk/yy2qvgvKK4dhXuA9sx9rj7TBghXqkbNt120h+/mDIbACGw5d
5DrRY+nmeXzRKW7UotZEg72i7JkmZEjFyqThSIyTb6kHY3tiMWhmSfrnq3jGR9oriKioodWadOne
7i9WEtdScL2+eoesX+WRPN95yWiyxUEpKxfuD2dzJ66PVBpLhzvOpukpo/gDJqNuPgvr3FETTtz0
vFbL7Bozg8ayI3sI4B6ZAA5MfagPYpH1CNpAGwzQQkb2Jd/f8e3RM5mK4kwR2Z1EHxCBUzPlYXdi
6T56f63yIh2MGKhbc4xzNwLt60ttVYbAWgmBf6PyKONvZLpgxhh5DD9TD5b8Dqi/kvmS0yCbKoMJ
C98CnttHzQ3vKkMidTKAVbfmW1rnDdH8iIpRC+nR4ZhFcLylB2Vrgx14L/ix3GAZVMQ8o/0Ta09P
HMbhINCvATRNJjpVEaZ4iGSO4+GFx6+1PVTC8dQCpVOhorOnu+patKHdytqtzGR6KvCsdeSKO9nm
QAxRrlm3V78WeIoWT95bSteViQWZjzG9rxzoLb9TIby1AynavTiDBwxqbHY80IJOZbNpVUKZffo5
ROGY0jIuTFnlxAQiZsnI0sHgA1gn02Zk8O7DuOZhfyZ3NB9jS0ieQIFQGEDU0VDyvdCK7OLOlVmU
o2zKzGKxXnFFLufJj4krgtW6Yrv1IuRPYkwfnsPzXM2WJV6359k14Bxg9i0Wbt/macRVDMotmYjt
Iu2jaFuzFRNa2oK8Z9FWQ5B/YRTAZsqaOvqvjNgR4q95ByuCcydOouEXGrlHQE+MEhYvIWvMaWq+
ktZhWN+/A5jPmFXSciD2aK25MM0z4HWItf3Lz76o+HPKvBlBCZEKhtBzMPbUmlCLRBUvzsUZNoft
EVyoR4INjnBRwYQKlPYugDuZRPUDZ7XZDl66b8Hwdmag7NzjphSuYeXjUVIAVV8KDGo5qpfJQamt
TV7xpD5yvcUkjhkCksGSGSRBTBqYXAnnHj1bLQf6VETYkWZWBKhXaEifTPfUnd2p0MtThmE7iqjM
+OA0Fx2y8iyRsuoHPU/ZV5tdpYRysmJZlK1PgAo4/HgTrNp2mkTRTP2DQSjPE+4Wl7anbhTxS+T6
uDI///p41Us/EzrxRpWAB8Pocg0FSqIcl1Xx4PN6vvxWwR+DDEsRK9Z0yLGJ4m8pFNCt+xuUsMHZ
omHUynGiZd73mHi01YS9A5ffnrxNBPED8eXDTLtVnDSVW3Ql9HH71uwh7X5wPZMRImKEuAY8onAe
pxRktTl1aU2hPl41s0Tw7RwaHQIlfgOh0sllmvjJUC8qHENMd6KAqDZuSMpIpR4WUDkDoG17m46F
ySnXzUB2JlpLurjapvr2HEIIEDKpDdmW7GYPQdQWa9MxoIEMdp2PnYYQV85OM20suzGu+ixiScM4
VPUCGCFXsx98PNh9J/A0tdMYU7Lf++nGS6Z6HAT4SohT9DoOsTJ82bbS4a4PNFeTloeFunp996zc
6cXAkteKLCaQmsGtb+PxUEeI7YaUyXMBDmL0mBUCgMP6EXvfc+Z8aSEFkNcg/+0rw0WBGA9j7dZp
zgJd9RzoBwTZ9PLXrm+0ByoJMrBIuXyYHaYRq5ABieJMHfsoQcl08pvAj7BsEL5in0GUk5FCMIqt
dxis0/UTzIBvdaywT/BLPCGoX4uiBuHkeakiIy3JeAI93oD2FYxwjon7yAmteohn67/MtHdpvYoI
GawSmX4JaIJPPKHNNJrRC3MCRse3mDTyv7RV1Wvd+AF0X8LNJSitb5qRLVUiNnTIeQOqdyEI49pp
urM/ENX54r0A/eejACyR3DxRO41bN3lRGUYxrhMYi64xMQL7FiPAwIH0F+SUIgV23agz70oLdUPy
iNlBAe6mz0iXtLJLL/C6vovFBRaAVuj5uCqoIg/An/R7eRTVqoaJ4VivJEJx+joZwqGBYkNl3uYi
kNzQqMP1esuI8rRYcyrQZe/ZWmI8xPsellG0YZBoR1lrdGVMVsrmJxMb2C1kp2OYb6O3ch2s3EbD
2Q91UGEn7iYq/2bI6Cm0LePZj8LOUikUYk1K0HKScS6Jg089EoggsDAMSd1MiNWMTpfa3YxCqXCk
BeqP1lXUCc3YeRAwIkB2kyEFUk6QqZYzPgM45KZK7nGjT6V4ElUnGWuODKITKOx69SbX9DtwNNdD
5jq9ItQ2iX7vpXMtKB16OUzKoyKnu/grM+qeHgZrG4YhSbTyoymT0XK2dmNtuQA/9QThBVcdGIOm
cLSAsXHCm1aqGaDjQYkT8hFdqsK+/QSICkScEpzBJuAz1Eh/SMFeW60MS3rgsbzoZLa4Edshke4i
XWNJkTJlkqYySRpEY0XmG+/i7AHCCbaK8xnJea37/DgfW4n6/LZyAi6PfBCmBwDNP8Ibs8WVAt2s
ZKUDkGRnFOsMqjinAg6kwNC0Inor5XbtCKCL9QYdIKk+5si9XuBfA+seeKrDH5dPuzRVJYhnU7a2
++ylenZ3cofPOtxu5V4OhyLM1AM0ww+sUG7qnBOKn/JGpcMyELs+kkjBjA6t7TRW6tQWEB+xdE43
uoLNzIhtj24TjH2YPFAUyP3c03Yat1wW+OYdm50EepBijF1NQvFLV1TyW5kP8ctuLe8fi2oEZOwp
uhwdffNxyokbMCUufjSdX3RHgkW60GiMQW+Gw2KYRrQqaAJXwMljy1g8XUKXdHP+C95bROHlMX0x
U71mg8tdIP0BgptaeIykfWxF+QpTjAZj+6zQVdPjDhEt8K53ZAUEqJ2poDQdnXuRCXh4x6xSw+uy
KceuO/3c36hExB4UHbgwCGk0KnLRySvnvCaI7O2cooATYYaNbXHzpvlsMQneh6qdyRreGOSAtR2v
7HJto+isfmRyk58pD/N3Sk9t6IjlsmpYE4zHub24QQbGyrXGq2p3IeExZ03daPYdl6iRJgbdzcGl
Sm9aZ91vQaGRadppGM1OUB7DF0FOce7gi6nq/X8YVAA7w6d9lA/5PKA2x+wyERXRWppeWf00eupF
gpv5j0xaTCMoDCVGKqLC/8XSbJ5ibR/j8Z+jb2G+kRUFNFnqT2rf3UYxr1x9F4oSPLhnwkcedQJC
Bt1UYNGOJC6NRZgMYNM/YJSXTDcuoSV4qy5ZVohGv3EyNpJit4gpI8TqE7/x7BA73TiysE0c2PwI
pakScAxLICaSY46+juUWyK7SqFdlIeemQWcZ7h3MiLeqEs7dPNjnCe6HLtA2D3OBF1iFTg20ikZS
Msst9+6n/s1kM7Z9a6unYANVMj069YDIYLq+9Zm3XxnYjssu4mCp+rK4kPy6uPx2DkchrLs00QkH
PZBbqrjESClvvmUhKmFJ9C7brSfnrv05lddRKUjWE/OdUKqjnjiVlkhf2K5xSg5NJZZWUOP52G8U
nJcp1Tmmxf8NdIFjm+3QVcl8903Likw45de57ufPXsKcz9ozwDCyHQ1xt1KPcN8krEM42ixPgTZB
2oTX00ARc7pAGFIjA1B27PUK7DykdmUayDcTIGARG4JgQCgUIL7xxK4hGc1CSbmbIpslPOTEF6vo
VxehFXwJ1h3vcSvJ7EixyXqcuYDZXGrXTZ8b8vEuite5nStXLO5/jpXs8Er6vkMskW/gQmumRnBR
6f8B3epCna3iBxBIx/lMXMcUCss8G6z3dy2swkZM9oQJxWDG/PixYjKb77UNd+w/rqRTCYr8Co1N
Wb/2EQQ/PePt3lLNLUWKthSEXulFQQ20g+zAQEGFwbwpD5luwAmJ7dXtwrHt7T1SYZJqXcjnsswD
10jex2EXPEAegyaRIcZB2fR/gi8WhiqZnaLGjS6B+9NYWjMcoPd3qBoC9ENahI4CQZKANbTnzvY3
hMuzH/W2dKXXJts6803S3uUsjR6vbxoiC/d9880aSYKdwZJHXjCxqnWw20PmDmnLLHLppJDeSEeE
4+1sw+g0TM0xcwvEHj3gjZc+glMmPO5yPkscst5C4WO6xOIYpPKS4M9/BzUVPSGNcpV83sDYUdr+
HxPPRzNU78ve+eGY84Tif3F8lZdSeEG0wHYlxwelZGaFd+MuqBvkf1ajuAhXIALgpTCxzkH3CE95
ASjyKFT561VHNhqgtUSR5yJETJALA7RHr1+CqOUowCTjvzo0Fk/k68xndE+uwaFnoMuc4QbTF9MR
ufMWRmNwGm0JRnlyPEt1LJGRYkCBsG7x0W+UINsfJSlm+3LsDB076lCkEjc7UETBMTsCuyaeav+f
AHzTNen5XZs7NVqWJu43OKmhvHH6BIKsZM0dBmTTnIcPmy+lWAW/m4aSZK/sGSwc+xwSocxk6BUI
IU7WYeMpy65J0GlbEyDjldIVY9iStNB6Hc4tEEIVYaoWiF/L1UdQSNzu3jLgK/D3qmClPhROLqeI
QSa8IFLIxfbKYn0/3wjhzRSTwVhqdfJSUa6acW7MyQA8nXFsMetRMNboePnxbYKFurA/qaShg8PC
OIPdEdgO3gUhyLpPcxQHAEwB55xKsDjLvButI+gzZRI2wSBU4KW78yUwCa2K7fWYFRmBwHxKMs5h
RxHgo2XTrs+0+hMPn4HMMRJlq94eXsnMuLwcBgzNX60FmUbspjW/4x+/8rC2OvcRNoXEyaU+3/SX
f63pjQ2pFWJ+QXdaHhWoTU6jR9nMHk7jKZhbFSFqCD40J6q8SbWrFw0OSsRN1jKhCYRFibdODeOw
Sm/P87iP1rjtcHCh1XOIUTOICfjQ1fieeK3fS7ofZ5xLXTkhIWIFFptd7lh4M4B7UzLHFAxj0KjX
eVqOV+hHxhz98rRV70yI8nnfnNyAcjeQ3doOKGE1d3mpZeFtVfZyDuCszCjhwCDTjJri4l9+kb3w
lpIAgHcFMQvIy98tbglaWPRwvMr2Ro6adxyuVxCTe8s+jKoJVLgGsrJaRM/Dhei5rXTMv9OSWc+g
8YQvYJSkGGQJju16qDcMNWkU9TbwrpCYX/pGdJafPK2s6t+JzXV9tuR5+69gGcZ2c70T509gKtjf
foPbjm8R7Ecv+Zp0fQY0ZcFi08IEa3EJeweoQU8EhzXO1rbaOkwV4mqNwPygAW3vpYjl9fkPv/EQ
9N8W0OL0+/7bMdR2STBEmnYgXzUauSuTbxfygTq4r3AGI26fQghCFdm43sXRYnlqJz0HTYrGPXS0
N2y1g5bUAfBv/otH6wfgPAghyj0DWWm4i6kCv934QMAR3Ol+RoPS+F1emwZvvfnoRMRTCZ8Po3Af
7q0RpEVgmoqCMXgMrhwJoAB9EgGGOVbbNg1zyiW/EX+EOeE3Jyy696tbTaO9nZSAKO9HML42KsEh
ckSgOHCf0U8aUISwhzrR8LKoTv8clLbezXROCHM/zSWmzCqXqJKHEKudfmqCyE1dj69Yx8EzDMOr
Eju0megvWeNlZ0YvcnL96+hzL8tG7DsZ63sGQPwwdBz8FvmYgedN8X9OptsJLFSb5RMxiCnMd7kQ
1RbTdkb3HU8NZHuemclxtZcsEnHuyRLOCxXelOkVSc+v98wfFUvlhBX2mkpIuaToMTONkrrDXN1R
Z2S/yzwN79YiCZjjyRazejW4dxKOFXwoUell3DiBImvTDH0dTKrTy088XMcSLxsFytYK9QM4/U3n
Ra81nEFIafvU+OgJMjkO+n5SvHWXsEbQLtVIsGxnMA/2+s73WCo7YdOWP+6mzcFU51s/pb0y/XlF
gFdYlHf90eEYolrenlau7Rq59HPaXFxYhYsN9JAIPy4OjtF0GLaBm5Q331HawBUhzrq3/3/5WWv3
RLc2xn5wzuLaXUF8JFlKbEyFnopfjwrBQFcR0rIPxAU2ryVII9xPmqPye1T+iWoG1PPE/6OUkCuu
T9CAAjj7EkoY0BZlR24zmYducyLVMxUK71Bv0mA+mJQlCjykMOA7WXCiSHGp0m8KJSYJkyr3N6Pc
fcrG/IZxH4iv/pVT0dXi/wm2SSs80hrgWrS6+cPA7Dyb9IARwNCYIErVVc1SVoGzwl91PY2fcQhV
aPSeOznXw6ZcJHps4MUNkGLCP80jVzhFuUn6/aq/ni/dS6Ko82J6ncl1+zdRt4DD3NNAoClhMFEG
B87t456WtIK/woKx9Bq/CeMDJynjydi5W1RbeDVTLhQ+bV+H3ejpoB2illLDgEpnXZxIGU3L4eUc
R0Bx8B/ZuAUxxg2Zu1G489f3Nbe5Bz8y3/jA7Qw8ExfK/JB8Ckg9r2+7Y98r8/tqjKyIK3CcTH49
c5PruJu5oZgRmCg70JtvUHbrnz3a+gPmJJmt8aRQZ7dIxWMvpVVeBI7kDCTBZEmif6MvwMAmPzU1
+xE9vaA7y1N0L6dXZFDa3LVPDuS7UxYkbiluN7ZUQ+9Ix7Pw/Qg9Rn2HU7PvHENj3t+7oHxwI+9J
B9fCbRYsUytTV9pQZlP6dbpJ9WFp6WeNiKCYoIbVRvc0pScLh+/zbqPIIgpgKdMW3OJG1vFcxIVU
WS1jdO+1WFdzIq6WpR0hl8AXWw4FbWUe2RhgMncpVeNoUStdDDM10xH2L/0vkKkbKT8MfIRGgpkr
cqyfwAlL6NFJWiIF47hAHifWj6/f+hdm8q6E6qfFHT+HaoUfxmoN6cmI3es/roHm7ukCSDrMfi21
rMj3OE9QI0wn4e3oUSwAS7GgVlLDy6acYvtcagnPZggpHPzR9VjZiH6/Otq8HTKXdou8Jo6KpFca
8FUaSdWqdrIT6fKrb7XG6C2BXflcvrgIGTg8T6PquxSeSwiLtHcmLr7n/cQ9mSO4GVXBEcnoBgjd
qDpQX46hAe57fm4pE6d/h+TrNB8G5B3OFUe1WcRHBbQ3Fpj4EaFO0lnNJuvFHgA7e9csQWjKDAqy
iPpUFpMrrpwjIwOIiZg/50e6Rj0DENC7JFzYz48lZ/zrTS98MGPuhSg0RVcmCx4aeJ296y2idWIs
OVik1w0lW/XL+JhquH3s1Ohsq+hy2VvBs44tYJIXGASn6tVJBKv/5A7W0LL7sirr8L31aUDspxpf
TEDNtUdzwR2jw2SM9Ghb6Jjt4lEoDxuXDTsBFFf0dVBNczq+U4tLWjC7f9dCkhm4roAaMI3k+EWG
tT7QTgeTLqW7zu6+Ppfvf4i/gtPZXRAKPMkobLx9vs7DOhLfaTOfBGPr4aWpXyJfE93ZGI/8UoHd
U016MjQIpBPypl+caCpk92JUa1jCmALuvzynMm5FuMDgKCo+ws7PdRxt/G3ABGsa4m6akCDu1bGh
wz5OkWRTEYNywSRNrbVaw08kLlXaMTRCKElpyyCig1zvGThF6W9SzZEUy/dfcoEClYoy9dDGlm2G
ojL1WuG+sUoFPgag2byelXrb/nS3VX03p+bQW8ewdlFv3LRCGsUtibyIsrqcziFbXRfcKAQZQA1t
yXR/JX/TETJ5JxeM+DYMEcM/xUnla66BqS82kEdTsBVszvfLPvG6Zjtlj+YKsyEa4qY9MYEPurfW
s6P72UbyDOIPcZID0fIgdlaFWyTUT7glNaExVsrsmmzsQcJKF3Sd1MwIgHtmOe9YEVL5DIqazUbC
TuDxW9ZCUIYiaCzVQhZhh1XqdI7ybYLZ9Y+TwAEV990cWu1nDY5HywmVXoLyM9xsqHj4c3bifDkA
ZIdEYvwip7FzMYbG8eu+fTxoH1jIWTCwLVad0CKsvkQUJt+vNDB0MWrubB9V7oI2U9kp3h026OGn
/O+YCM9hN42ID+eLzk+Rc5IaAYnCSDrZ7v9f2IyZUPDfJKxuPkaBuccIWuvafcyFQDsdA/5XEkiU
FkZmGta7HRdnRXY6AjyEF+jKV0TO6KGm9WT71hhbwZgUa7wLyNLBFWGzLFAgdIqfGkUlwQQ5j/7K
sBqRywKSUK/lOyliZMmzhCAz8sDQSIDqMjyv90OU9o9a3nkA6eF+5Qp6inX1SgS3Ub+U5qiUeYLh
izRwodM8bwnDTtkZXhUKUo2HlHY25w6FaiWd6uD53SiX5MW89mAvye4cpKSK6XNnwCdxKPRmrf1Q
YdcQ/0zqgWoQR2mWCeM5OfbdnDxYzzk8v0XaYGRBcc8ZJhaRy4o/gnjoxnypPjPVQqro8xMUBw/2
KNYFmvgepQquUjmyW/tMQGot7PVA6eQj9zO+WZBGWRQxhDdWtqhFPxee0wgDvTYvjIj8VxZn4EM1
hePybjapfEPRWIV1Y/DxrJxojLDK2e+FxYLGKhe2bBYhvbwhT9709PLz7UtsALcOkLXEFW7oYdNd
FPnigJYzFeWv586JTOJsoTrEenE3OL12T30BacEwEWcEoc+WLJsAryYgKxOuCPhwexUbLWAXj9fU
FOBSJd+hjl6LMkPwnFNrjBv3Nuaopk+P/kkySLlXacO2dZ5tFcfL88dzzn6e74XyI0Nm5pM7Ytiz
vzs7vuyVozui6WXV4Vv8NqP0k4ONOFaO4pE3uEaRG2ST4lrECq3EGaY/84D3eoswuK9GAhIQ5Il5
UhS24P1kAMV7C9LkkZdMXJv4wTWqJe/MwXhoZrPv4cPhyGJqdkxSrftbRbuwj9dgpzghE0s78pzI
eAfjCj+eNi8KTi6rh8g0wHiNjJH3vENQQQ+ZTm7eV+TEp2pgnbfKwLKVMtEQFBultocxMEhlcWvu
R40ijce0HKf2/vr1oNqzzIL/BJpz7aDUt6zo0QrUR56lBe1IQaTeS2Ja1mf2lyFL/d2hG08k8uSv
TnLRaE7WpWtHbnhRYrGnXReGA+tlmjyOOE/+IeN+40xCUwnuUXxui5MUo4/8FuNcsnduow3keMjw
E5cWaAYUgtJlh47wbe/aToEKXVeAMYffIvzuG86BVPbKitwDaU/y4DB8Wr4rSP+ZUSfo394lP01B
IibFCi1qtApDtk1kQjWJlYquy1p2DenWEIim1tA2tNsaZ5L/QqRyAcbJL83Z1EkuLmAR9Pnm/uvE
7vSI1oAWFPlUHp6IVZj/59zyUXVplJI2ZNMbGR9EJiW0l0g24aQXIE4NvjrECJ1UoRjQsYKB4+yd
jXQk5USCU/bTDnEOkXc24wad8/2FrtknWRKiXj5lsWWtCbMEkhIFZ3ldf3xbwPCcHsLT4WqBcuOA
vi0gPfPX+CFkUkEeU6w70TBsTmaFvsDaxbOdtHirz81wJi+9m75k44ZCP7O1/ssv7nOT6mwuBZ66
9sguADENOA9ZVCBEZvre4oUfAGYQ4hEL9e99DrZCs6u0JrYaFH21nX+I59yboG3UQtAbZwM6EyBM
JknZSN0TG7R9Qf1MN4sCm/jtM1FENQQRUQCx3Ef56oyPZow8kR+SDtSn6qFrAu1Fn7QEdPJoW/WH
qv//xH5+Aagp19TTN6Y2ARDw4KhOHP6KQnk8TIVTbDKdC0stka04ezPvmntpXvgx3tQGgPLM5gnj
tTBLBd/bzw3pw4IPAzXwPT/jEGQoadhOWLOnnjSYyMWBddKChgRca2Y0+UDVNciDeGmevnX3Q/oD
COgpFfrxK2MCRz/SgZg+AYyuyKLdXQirBAvbxHW5vqu33gP9FiDy7lu1nHbAHULK3IOVl3r3estJ
n6Fb0Cre5OTgbhhaU9ex7CRC3QtQZHTg1EnUoAbfbsEMPvaW4RzrzVsinU8uMC+wSgIwNO7Btql8
uO4nO37Nx0qsMS/mS4LUV3msQMOaXNO8euyDPEJQOjgj3Bzkg+7ZuZ0C9e8yYLtcfHhffxXs8Xt7
xrHLw540o2GlASOvV9MGF02V4DxnDViMqzpG3g38oLLww03QQOJg8Dw3kcl0q+7D37PnWVHfvm9D
TeoOC06zBroC+nZxCaLxae2EAtoqK6VuE7YZ07bJsrk0JMYEp5zmOXcPTESi4HIYv5ilhsVq92U6
+Un3vBaETXtXA6DFmN4/V7OAKck+MAJqTpHi7gUFhM9m3vKYkudmtkRxZsBIhpKoBxbza2IRPDBz
LI0jvsPqhAIu6R+OhTI7NFnqnUoZ1960uqL43jHztlkqFL0IOT/tqJxa4BvSSutM7SHnMPjfF+8/
JVovd/X+oSXarKj3kYDKzP0VC7TG1JD7LTcRcwvIBpBotQkYcuUQIXD39c6WIT+ndE5oHcC9YLAJ
6oX1hc3gJKiz3XuyZuPY8jA/490ZXwehwV3jJFbFJDbdNEonjR54xclZkdxMKspef7Uh5uMn279H
gLACIz83DVwZpYGpD7UnV971+hSRRSt5zDPAM4w8Nqn2VDRj30b/Quydm+PwWsyyxo/PpCASuFOM
8vHAayQrRA3MwyZzVOvc4VU6nUUkiaBQ6v6LnpzI9kpz8419IA0dJBl1Dcdrb6Ccgl9/nkAIeyiF
EHQPhXtARP5NHccZ2NsNeaNJmRkWwAO23l5O4vKlDtt1aCKywHWKLnD09E67NaVypwyXap52HVuL
8LvGRZ+BCWUWD1PEgZppYONglRygGCHovGDHoCn5NlbDqzCt0G9oSFPS7IEFWoBr9wj/7Aopr+cT
pg2AHNUO0KBl+BTpVvGPgJIrOirZd8uLOcg9p6lk8PquszRVQ5v9P6ShaIAuab2nKxRDdqC3+nWt
Rp0UQLPg9ymT2YgoNRCdCiYDXklkagEwfQpeXuuNhv8qkeJImKfGvgrOTyVGI2Q4sdp++8fzP7HI
RHWSlFQLj8I4+LfkWJDVAht425S7Hruv9gn9Lape6KPL6L1mom5TWYMtGjhTVldcReUdN/EQcjvV
Y7E96t9IO2wT3wsYPEOu7xfyqDP8zfEYa1H4MwDc6ttEvJcTC0+GzGPirx9kvSmXw/wfaQIN3O+Y
hq7QdTXZ7pCdYaAaaoCFc6U5YE4FEFDfM7I+wUND1yhwGDHgQV9nGLs2PEUr2RFhskKH3kAezjFZ
3TTqhV9FzZUdF+TY/1sLak92SLb8EFZG3rJOSWSdu6MUrR7GY/DWmhnvDxB1fVeKITaXOJClxFDZ
lOZj3h6ilMAM0D3Bww07gJzXBwhw6nuHv02s+saCi17FHVrZmc4U/unEMVhuHM3p/AexwHgQpF5S
srGZVbagsg/W5Z0AaA+1dS3nlsTBqft/Et7AeYuOpbxwNTfzLyzNW7mdPvlaGo9KWLpcVwPD4SJ+
ZB7MWFMBrRcH5ekbDPSyJWsC3FqsaU3u3iFvj+xEhqibzdS9E8T7ifvFJv+B2DNCYVOODNi5WFOy
dNU+iBCLctj+WWBo8k0CDZ/6LS1Z5aOqwdu5b+jUwd1SrVCzrQBWpUUxAArcbtiSOj/715e2jkDt
KtJRAuIH9ztr3t9YrDAkoQmPEIH8pA+68Mhks0meIo3LR2DZg96a2cSBNXPGCRmOQtojFj0sEHqE
XSwHdSUjrNk4EqDuNbgbjFvUuosIjQolTtLmFuuovK/7+j2XzIJ8sp8sFqnNd4RvEvmWj1ageO65
MrsZBl/iH87u0lHbkQjdSkfpknpBV2S+wx8JFouw+ta4iAhWJ9jm72tulHtY+yNRy6CufpE9wWXj
eY1X48KdcZT/a4R0+DhGeZlV/aQvW8zbA4crYScvdEwJ9ZX9BuueYko0lcftjNd3HOcDRLvAKlvF
E9P5PsqRg/C9VHt8uztFBbQyHiQlLG/0FeylWdoja2Pj5+a6ArSn6XFQpDay92J+I42tgYAMpMbS
KtwXhgWTiOe5WI2Q8TLeA7qPGNrEsS+aCsroDe+ARV/Pc9Yix8YFMf9KZsLR5trWgjDcLsgj2pyQ
BA1mBJ3rA/noOOC4FWnnr7N8ISE6JptKvg0vpgjs5vNgecRHdkoeFRkKt22mVKiTdYkXmkn+53M1
9hUKCTfmuR7yLeEMwnOkvXcBmudCXXrh/ED0aImGGBIryrP9J/IapxA0/HXesGvlkvXWmB/zckBt
o4/ktO+mvDTunmjMGd5nddHJTUAZaZkYAAjsOY3wA5PE8VZK2g5qfCxoSw1dDu3tKdQcHksEgx4Y
ySUgCQ3K58XFWXkvn0aQ7P2WZ+W/VcrV7S+gRNpNe7OrDZh1oME8wxSjjaRvhI/N4Yj8jyDH/eKk
h8gMtogesVenX/LCyvm8PMnB+QcAUo8iYhrKTHMRyKR3Fs/MoT85SYnMWbee1wKQgCv8E9vrekty
yy+Sh5FFZ7nkqZW+L+6Qyvp/M2Yv22Pi3TwulqTq9KCG1NYGUznHZST9m6qmjXluzcCzlBVKksTp
rd9rRJ5cv3QFxa0NZGs3BJtXpVnKLtUagK4Kk2WIqj4aoE1FZeEe5H2QZQfAaIlpKfk09OJYRaVA
U3HyFPMYyNsBIv9I9JEYi/qkZh8mLHh9cd6MWefiIv3OZpahQSIIiXLfclVb7DbZVPBQdsm13Mif
FpJV1LyEc845pEPxgWM28cVUQCZ24AaVi48q3SE+BiA7EPGQOCauqZKdLaWuFWo9QqOGoOUOW3yO
F14qDrNOuXfyuSrvd++fQl4ZPuC4CZ6XkAI2iMw1NSWE4E28McGEUvcoyKnD8G/OE5Dq4YSWGo4J
YioU9bip42A8g9F1IJX8ey2fmAHVGWRBNX9rH9CjNCYWsJLiCz9TVC+nnpjX6zH17XUjPogpwVP7
oG+bhJ5tuaYFFSclPt+5GMO8BmjrFe6MeGKKK+1AQ3pCAXNjj8vL9RRGTF5aZRfZO2UkxJm4N61I
9saJxdNmVL4Iy4nRJAGh/KJlnl/tKU4poxM/rgwRrwXaUiaQwN9V/Ayk0hhdGWNDYcCHXQ7VRhcz
EafG4Qssn8QqH6EL0j/OXWAKJOiGwijgnd6X0vO+r/j8HQkTtCpa0TQfsnccfUIC872bY9QwnQDT
BRZWsRA3egR1EcRlRBvwevVUKkaQzw7UEPkBxTwxaBpKfvkuCwnjhJde8ZpvaNYg4XRv6jZcedkG
dkt2QGlLTtZwaiqeI6uR8gnMiFSXckIIVHi6bYFGVc3NHMiiKYLztK6M9D87gk5lEFnPkx/Gjp9X
BATsN6WUrcHx2bYjiLJhK9NTIpieH/phxpdPhCTa9g9DjSrKrY0bOUuc5yLgZvX8OyjmSNhw8tHJ
1ANGGy8CQ44mgAEm3RYKpfut5UB1aRvjXD+xFtO5FnoCWql4nCg/i2Gch9CItastvo/SPrKUUj34
X8wb+O/Dz3/sAia2tzXLuIjpb6VG+KiasDhIPYakDgvYM8exBhfEPUaxm/6UCeCjfN8uA3lo/vZ2
6IQd2IfcE3B4x602JCpjzqRH7gLpheEX/vBSbdgDaAt5fjNVEK994tijuLq7dDj7xhsiibO/tZ9l
QWiBbGdoa4XZCqaKSCkqE/4bP006QNZnQT3XuVHNXcs4/EvS6HQg0ERu47ZBl1fo6qfSXLfWWOGx
4LtPqZWoSU5tiiYubt9d/+vAHEE1lpB4t72sOLz6dM9VnetXhDEh5ElhxpbA/JondX/V+vvsgz9v
ODFsJAXEQ1GoowkCdKg/AfGdYO8XgX55qriIEUnAmkFsuQzNy+2MGgR+BJmAcYf9t55fT6+PkTvY
DpP8dSzz+JWw3b5b4JmPbziQUgi9KsakRXblFtajSGa9kTybaqP9/yClZdUEyDoA25bXICsM6ZYI
oMIZECnl6kVbOWy1ocxNw0ipqBo8yRBnUUeHicb8+9GfopPj1RPKBj0tUU8u+zEcnPmmAa8TLI6Q
E5ehk5LTrtZSF8/5StOHfvnIOMm2ZY+FLXDToSgSOPctCDw+Vv73TTx/mFWV5x+8BcAaFCsPcWin
Nwt7qDO9gLhECr54JvwetQbahRY6rrECgI/Zi4ROmkwRfkf7LZoUdKHitbPn60ll6YMkh5ilZ1rI
Sdgarw7OXxWFzH8kMHxyoI5bnLSrr/vCtcVpijMzeJJzIvG1tMC5HWcC4CTmuJM7nbIaxWGP/7hg
1EBTB12hon7dFQeBI6k6m/islYjY/J2tEKz3uLUOh2yh5RUv+nARwVb+qJ2HrVpxBtJkSSbuXLrq
Y2+xMoz0E7dYmej/an61fj/aHIw4JD3NwBwcMbV9b0GH6aN7SDRK2NBnrdCYchuza2JfCbIUWpc7
hPYDj0FghwzaGp7NmqpeXWtqllYSOAMIdbuuKXt/z2bw0vbCqvNphbrkHn+E1V+uVPog9THGA9Da
aSINhNKrlZ2ztxYiT45yi/EbZMPQhlaqJWND2DnYLLQgTtlZlIzS9TU1OtyGt5uaJjsRCi9dXzn5
UJCvx50xGRAIn4yb3qw8A3BRNZQa4mmZ0ATfxtbTEaUnJyTlHItNfXMUnlokwdZf6ouCjXTekwrc
cmfTw2l8L4Wr6mSWNdU2tqz2Om0JBSFmG3pvF2wp2UD1No1As46dqMNGdHUrIZY82wPUgNrHcl28
YIaqk2ZbYMwpbWKhPDdGXtwlGC6u9w/uzlwc6VXg8yJMre/2nZGZvMVuBXrK04mmeEMDEJhxOhMj
xP2A3fjYqao2H5Tdo7/E1hKsovvVQ3ukb8nDJ+RNnAIxs5V3MSGIWiAzDiyXfOqZYTq0N0B15LYA
2AjhSb4837D6TJCGSpQgWfVDaTehOQzerGiQ1reaqPHXTgibmB7GQl4hBS7iLMqdggbAR7xPtOOr
H1CXdJIFs8vPfLyufR4gRiyxHU9W8w7Zhyoks3Cg9tJLso2Ug7XSS1/iiuU4NPq3O8RSGbp4sx1K
cgmiKJJsiUWrKdEZWVdOOTM7puY5QjJDrMDcK6VgoFHJGFxFWQ6lzoKvDgEWpnJ0jv5tobDjheTd
d7q/AYBudokaX0yriTTTRZQx7aL5bU8KDVPQlExpMKkD/mIqbqSlhr7JRijHi077ctsrJOUUspTo
s9b3gDurEckHSVWeh235BPTE72nHhIDqRUfKPAzYJ7D430cLkMC9VzDwY28rvQIvCyN2U8ZcMgl6
pGN5OJMMqsUPPU2Ba1fPtCedk4E16ezefb5RHQ9uJNheyCDpl2WwHbGq6/8hy9aXzy2K1DRZmTlE
1IijF0xWMNj2E9o2AdfKxUpv7PDV6Ms+S9v9m6S5WzhrajERZJDm19ohrLzPE4419dHB+pFilQgt
L0zxCw3orqj78GSGaHAkrxbw/Xqx42DTZFA+dsmc7+9h9sblqTZppHBSNN9mJb6MKvEJBuPpcHFQ
1OuVJBPeHmwX0dOowOD7dREKGrUB1IxtTGRFTs51w6eoa89PwjWsAJeQU780KzYSp7D7WP/mDsZO
O48o8eAf2VZh6EXFw3sC/ZNe18VV7VuQI9sPjyMObEfbNTZsAzdM6RFwiYGvVQYp8pI5CYt0ChCV
F4DNjGXx40gUyYhS/bFNRY3t+TwBCvf9w2RDFe65jjMkx3EH7AARngHqHQoNZTigGwODbOg1gQHd
hn1pmTUorbPqSBFHm5shRWfjpxETCduMEUamTIRf/jJKgUxJn/Y2Wc4uCcY4/0ScUe0qGs7Qds5S
dplGNQ6B6hpcIBpyXtlMZljKsB9Cu3yPm8XsLq1zlDrw6cDTabMHElrP5q1h8Yjb8qNy9nnqXl3j
nBmptb54TJX9DadlGHfkAM1r4JtLE/SuM8bjqYnhbrmp3DffTILEn3Nf/4zyJuIvgTCR9b9hPBiS
HxraI4jz0uUimaOnDlk7q5FNe+6ZScyfu+oVLsjIRa78RYbfS9M7mqOIS8hpJDCO6ujCACUb05xy
phe6+Qrqv7zVGn+jxkFTWDoxcR6rp185aB4c7UttBYFBaLyccTqkAiGduEU40OjixKr44jb0Csuy
wwCUjCcOrP/fB2IhNBM/Pj4jEL9FXuzVmwgTUKDWtKvmr5qnFTXp3tw85nuTtsPGxveiJV2fYWWA
1kFrr4+zNXps7aiRyFqhvlHffwuouwbUOLSl3cw6zwutjSVpPELVvXsXXunOQ7S2kTiu18ZDFrU6
m9uYkf5HX2cxCFhfYyX/vYybJ9vSmX1X4woKq3PCfxE4rCJ+QiKlljuDa3kMrtdFuel2B8s7ynne
a7M/vFw6Pc/ZJqD8mQFFgsKJuMKIr9N2FOq9Usboz08EpAmW5UU4jXdqQgyXxuvtsVOoS88efWQA
wBhZy/JaY17+dDEWSqLdiCB5G4nKrt0PSecWrxPGwW/31WlQ3CI9i9kgluh9xmHCraPmlv+NkfKI
7q+OfY9vOh+GcfNdnDUaDAi2dGntCgHb2wO+2GMpKi0R9eV3qOSS2m1v0s3/AtLTrBKIBn9UNIY8
1mam4q8NOJ8T8lmVo0FPqbCk5Og02xBjb8ppZeFgjxSZVUVraHopBD9dyRodCnb1r9hEvoINAv6s
/Vb5DZOTm8yGvhuPUm6tJdjOHx9oxtALELxNdCJgSOkJqNro/Z9znvCdTJNoOFjOEJ3MSMBXuqx9
2xq73QoEKmSlWcQI4BRBi98hObVEjK6eTpUxu4+rJ+3qpxmeXckXEtJANK+4zlM7sQ6yE9lEQbfD
boo4df7PKJ3oKYglKV6ZX3bmgZjh5VbfJdY+Evvl5oDW8el+OPgZGtczAPuPafiHvkkIyWtZdy4+
1nHalggsUplP8E/ZM+/IMyRjSq3NfOWnJhh+rJj68didoHQGeH9WWwbnHwERH6KwwyUb/7/nGS48
H3gj9A+R5BMVT9VoqjCQ25D4jTnypkZIAYAwlglRDjgJCAOIypYaVesXyKQ8q5a1K2S3g49+ycLJ
zeU4mqx0I5T3YKTTx5PpUsL0gMWILXC3uwfS1GDM1lzIfatB+EHCv4MZidCPsU/ePIwrFpQjQczt
bGIcHoDE4ohGAsHcfbUbfmXta+/S7UlRj1lxYJO3G2LZGT/Hm2limzTRDvZd5cieaCCMkGYN122w
56rYQGw9nHwqR6Pk331YMgcXTSXB4xOPXAEBUq7k+/uzCQ1EB+iGfJfIe2gSOfmwXv7sg6YDAHx2
IB7eSiOX/wD0MOo/de5ts/ZFwI4XmCmYzWBAWfbYyb8FxrnlwdZKWGTqk4xbUiwNbj3kNYZ15Oq+
Qb7tsZRhWdBWqAuPl2gqhB9h2pNMytktEFOQgSIGYHFON598ZAuZ4cpqS3RJL7giCWkpJk6mcy4r
c1Bg+3EH44+K0R20klqvNHXTXy3BBxLCJOGP+AmZTQyhvAfblULDmfd9FLx6JBa9GoRbJ85zGTJf
fitcW9X7jFxSnRYvu2l1WwE/lPlHulg1UTrmA/xnEctRraTmCgLqqhtXiJke5nA7AJ9HKIUPWLKN
ocfKAPqjEMpVfYDnJ+dAbyzir12WPsrSnz0VYkrV6MgFWjTI0F6g+mb2EJJJVwxVI/5fy6xSL39G
iSYY3F8v9IuS4csST4ENa2PZc7twyxwsoNAmbJ4RGvqkq+PZlQSPla9zaB5FxP1uKutOWRC4R8Vr
h59hG/MqD4t0tPlqOSe9A1Y62hOsv/z8xDUqmaBsXOGKQX02jIKZRlzSFS403JyT3hZo8c2OdiUx
z9U1I7zPvKpcfv/x6LHTLDugyxLukFJp52aK6YVGaaJspcikncthOzWLzbuu4H+BHaM7HIKKVvrK
WapSt7xkZfeMXt9oHtB9zXlsSRI+kbuRQb3PkgASXvdwpG4/ntREGph2pKqqdIZTqRI4MI4+C4KM
VBziOD5tnEbAlx4Q7PNH0UE3u1GJqJcOAqkduibgyh8Nr95pjkQBt6/9j7tzGg4IrWqBCylO9Uqy
Ajj9ENvl/7tZtdSHVbeA/DNncm9tDR4BiyJtHeCdzNkUgN9t1mD6SNHi4ow3mnb8nvfi9w2XxTsy
067T3PMgZAbRO57t57E3nPflf6ywtk7Ye6NcJs3FDaIP3F7d5BX3IxLrSNNm3XkQ1aGKF5HdOg8s
Zj7Tpt2VtnfoX8kScDJ5OOI8Ml7uXA2DsXrZizQBmvhrZf/clMoMRxDbuHN1JBX9rMnSy47P7ObS
+onh8KNstcImjuQlQutKhMPmvRN69LatoGV6ea2/hLp1E7TgqoTChJ320pBvtgZfCDMokGtvmbe4
A3dudcj5Vo0SO2MfFMwVmqMcD6hAP3cPdUduip9N7V0xkUcdvo/PrQ/6YGrjqKcneEH96WpGk1R9
ji5cQopu1ooMP+3MoK4ZC+HJwEDqA94+8DLVXK0kdkRcdlFUcj0hOlxZqtc0pkbdSoxKPphk4VPp
7AuL3uHvxpnn5qEo5kL+IloGjnsc1cHhiTM1kHQ3inB2ROQ24+JPpsMpVlDxCqvUf4LZC06ZfzIr
HRUFTZBgEWXaEZz/Fi0XQvT2RrSvM1zlK0kwr9SebEOYVi7MJotZUCeO++zi6pSS0lS3z1C5PHoM
rHonjeoWgdeOntVwRNvowkApaJD3KOlIhr5Hk/D0BTAaJAF8sd5xoP3cwO+gA7H9TJ3e4COyHP+L
8U2D1tdbu3dfPzaSFUG4I+Ej7B8HjNj+xeRG0wT7/I9U3aiDj5KeuDTFvk9AfQHz1hWS5IiXA6sw
+CQzKFXT0bOq3ViRbisoFa5jC2U2K+6iz82fLyhVW9qKDcON4u2GKuEu1UPDWzdPUNo4oTfQnARB
YNchx7yTnl+EazpOd8ulec5c4U3uhVQsewa3DpU1F3SOW98+MHR4hGZ6VCDso+y0ODeGHfHaAE2i
eUvcbANQJqh4dSH6w11Myuk7SdbDLRm3t45SyYq9xtLEQC3rfdyOcjR0w78YnEgAZfOW+W4KPyji
FFKJlWOsMXNVeNg2Dk3XNf1b2vCwE0Vs0Xi1G+MDABafXm6Ekw4j69fcH54noHPvyAPjsldZ61Be
eRJjnCyR0K/XSUEvtEfqErNZUm6gpu0bKduj+SQF6WD6s+SAmqWCo+rUJiNFxDjdQnVDte47E/qW
uQXenMzC+vtMdePi8u1RT6C+3ZyKyfyn61C6NXwIHGzvRl5pL6Oz0ZQDMLNrVWGrx6KoHvOQkKSR
gcfkTTjpQW+/iEuuxkCDr8e6xVh9Nfqn6GfgV3+RXFojWhexTfUxtSNYCk10/xD2Po0avhMkfEZy
JcclM0zl4xr45A/vBfljy9eYKtPgQ1T7Z+ca9B9RiRpTtT8tAsX+u1eR/3fL9W8Ndg9CPDebQkxy
FqG51BcU7/qx1IL4EI+RBtkuQqZGihxYpmADhaL0vllYLCbJ404oYMxg4J1BcHWc9ih1wf8MmrQc
1kaD1+PayjrPi8onvoVV8lIQBuiLBowwGHyqBKmkLeO8WGV7DZE/EELUIAZ9C7Z2uK2Lrwv3VWlg
oQHsggFHHzpJKrnzi3HE22GRv2J99HsQf65rLkAzyc7/Z7ppRjIA5Qtoza+pceLB8MjlGEWsrjWt
sNIdtaxbRvm9BBfCaK8VxoJwWk0IehsEDEbynbGeQ4o2mBJPAgCcRA4igzIbLuhLKSXgbhQ6v/5d
PRxK6Wj9n3SjKfwAziPozvZe4YKI4ooo0HK2hbuljedfIYKgEbCd6IVtoTzUkslLNFDlQLxsYTz8
hK2+I24eMB5OS3cHL/XgJpniB5h56iflVWZQY+j94EGtDh9c5jSSyS4c6fhgxNAL0MAEIw65vIzt
sNgMYb0ZapUsSwUPTu+1tUNv4EcOKgnRZs1cUIObZPVW5vRFwXPs+ycWkvOnVb5TbDn7bXwAjVUw
udREbq2WDvJ1hOjzRsVGw5MLCcPpGjxVkK9sBHf9gqEFwLpRC2aAg4tFjaQms8+q9niqbWiUIQJo
XswtuzUA4+FB64ldMAOeH1EYQD197raBO04zkxSnwvQrI5DpWTdrhFikZPDavIY6iE0hfG05ry6/
tIOCRtr4lQ75d1BVuYHtCEIYeHC0FYZjrdc75mg7KSWDwk41OaxdeF+OErF6dGIli+jtgiT5vUpG
rnlzgGybra8a6aCvRc2f/a6yf5SYS0mGd2ds6CtJ2e9k4UiYoxPtiwuB3bt0LnQo+Fn0YxfWKsGZ
R7/ZMBj0B4xCwkZnlfmoOE+g1OeYlCFoHL8Gw4pY7ap/611Pr4KNpPVRmlaJZnK9CuDOxrzBnmgf
/7a/eFsFvP+8qchv7VAqSjmT3UK89OcBZN+16h92//9dQ/jU9dyoe29Qm4D/imRa/Qbm5aBzu8s0
HfkHzKqAa4GiDFKNY+yN7inQCTgxrpjswBRaxnORJYyImcuCLQe4n8J3aDIZmlwSSyLtlKrFkxhx
p7/eAQ9q5tdg9L1qL3/phadwOEmfQgWXM8Rumv9HsGsWI/qpYl2H2cu3cB+vaOnwME4MxK8djQLx
/+OoQlO49ivkLCPDElJOyt9EDqJksjep2B06a1YkPecEVF8AMpDBsZPxLmrDVuJRxTtxgKofXrYm
1cOvH9Gk2+V5bWcWb2RPtqXCWH2iVapOPHSgjKtL0m1WJF32D1Fu7QLThxCFnxhhuS7gSdmODOCL
r0+c8NDXIuhrLoaGlO+0eCcXGCItWA93QPWx4zHAkRkO97hSnGlf69hxr3B0nwjFF0KZxMmS9l5x
Kwso4jDwh/wGgLk8LTz/LWBrCtxpZIZo0xLF0fYponxvI4LfD7CLredXgOY5ez07xK0jttVFXGOi
D+2A2Cm9BxSYf0tArgHjXGO8voQtvP6jh7XScTsadYfIeThN9b/Ba8sE7XykgFpfsiJLd/pJsSVw
rYyfagTQsSnGrBFkVgW3OhwkCuRvUU0UFQM8pyDWRLntEmlNO/LQ+vQPWb1yf5tDD6zyG6UhwJK/
hzDDmiPV3P7FgGi9PRXfgjQxl8jmgHlx6t00CP6O7m6MBlZsm7IbT/SZYCelIYt/PZ1HFjnbdt7Y
iL3TYlEgMtwFYHHtElwGUhZ254ZXEzPe9jzdSgGBpLq0uGwklfnXD5PcLCMFnhKi0E91eUQLqiwi
4209F71ED/38v4s/ePnv8LNlJIl5EkS+KA6TFOIQi5Rv49SgTFcuJxCwZXZ15bMgTvEHnQfTaQaK
7S4HGNUw1sHI9g+P8eodx/Jy6amFpfBxzuzoNg22Uwbk6F0Ut4foswaVa/3pcHoTE4nF4ofuOGaA
B3/JA2TJQLL8YaN/AgsvCBBGUHF/cRwhlU8Z0AGmiGmD9QrAWljsKeAQJLiKQCa4Jtv3b7JKDIu+
SbEY+TNg3lSrvAhGy95Eev+/PnWVyj4uaXyev/c8KG6Kj5vWjUdHBYt+SWK7v4aD1s3CmFDR5exT
AV2XlptUsV5MMLh28I4V9C6TdmyNuB94mgxR3S5b1webTPRtXuRrlG7aTCyWoido150aR7UmX+J1
lbz/50EcQrdfi3ek9y3puowt/UCnOQrhlUdx8YzhaSru96r4/9yYS4C/yllKoWfUMDZt9+OE6/ne
ZOo9l2vXb0WHqMrXMRPhpMoHB419PIW7kXL2IhGlrA7hqZPOflVcUeP+4GaKwOtLwz8keyfZGxLs
NcJmDEFleTtmW3v7zp8y+Vhv3yK3Wo7T3u2TRMI97NnElxewVFukstVKxZgs8c+zU6yy7E1U2pob
3ieIzZM5PnNvzKnRoxXs69ZrMA5jYzJ3wSDMUtCusaSczegDtam8AyWr1/DfIAvIV9qHzeExhqrW
do/8UpuHHOl6VqwBjc3kqwCcjJSjmBH5TeI3H82+76HUPIoOnAvlwhH1OJWGQbjtu7HI8bJYEUTt
Nd03+mrTAbnngtZPdvU0H+CuIgfqNdkvg8r+4f+ShI/FFYNTYpC7TaEi8WwgsClBtPE0YIYawtsn
wQyF2lpqwn5coRgJsZuJpeyDjhXALR2d5dA+o8a92ZOwT0q1+d1tSnpMGPwyasUkFjZXfZza2Wtf
9lrSgPEXYt5xxoD3RpKuvitdsZI5dETwb4ygYuDRYxIsjd04HSPUTS83LvNFU54yq2md3ipigGl2
rakziCdQw15wcBfA1ukRYS2IuYXZvu1RhtNECiTai+L1lnwr5y2NhQ9apXjhB3Z9whRuSs7/X113
CtYO6Lh4gEWLPoUy7eI4ZXBbDWrYc3Co5f3NLdHYrdoDWaaRf+maaPQS9RVeLhOQuIQZJMPD8JyX
geemBV084G+W7rKWgUBKQ2zeZye39Tr/29Ug4QCnbEryb8JSoECy95CLgp9CZsqIH8Jhxr2Q/ZEF
4sHMopfSoaKKrig67+DQM4ADC85t+pze/mCVPfW893HjyVylOCeeyYOwb03yXuJ/KOAYm3Mg7YMp
jDYEp6BO18n+tVfgSuyIgNq+HGTPZHDcz+uo5vO1s7T7q9NtpkVdZoXqeQ39mNiDc26eT3YzOAI6
zRbNDuAAs7xOWB3C8kK0FqF8Njkuh/gCTzgZlbxkhn7OnQ5Yw3Ope1Ue5guxf0uGeFZPt0SEKOBA
YCMvsOK/ExJJm//BxM8GhhFSecQ1tPE8/gjVnfK21q8z0Aj12kgmywSycRzC4+MtBnlMNVx8qOXN
kQ9Z9e4MtBzwyaBQLi8JzbCRrByy596IfhQ/s1ywghR3CWPDgyZfprkYrUphje2UFUHBBKFinaxF
zy1/D5u2O9F6bpg21WnBnrSL54rFnscWFscyDjMexAFQOnPHFN3S+2fyXhcziATPd3F16EeNqFxL
6l0E4+6s59UofU+LYRCtAxnOhvNDYI46iKnlNETPpmtfA3lroMr0bA889d43AUjru8eckwxxI+zL
+gSlGYxzVjrMvhIOHAzXTS2csjtU14hKDlWyd/lG+geWzCNGZjjS/hobNF69WqfuFnGTg4pMqA8m
G8eUIm+QG6bcsuW8btXBflKLJGSPlUyz9WYxbQOpdOspkkk0exKwqQMlV3kPZG0qfR1lqxS+Yo/L
FuvE3CpKPtl/+Vh2cc1ohqxyaU40MkeasXYGSynpOfVUYOFA25ZFErO0nC708/+kzcmsHaj8sHFR
/SZI7X8ie8chXOW0mmB69CEYmSip/2D0x/jr6/55scZUm+IslFsRYaTZeXVesTBULGMMDG5vQQiB
ydqC0xn4pRQJgP+RMK5Mcs6jKqI3M1rMulY4xvvxr4EAb0YPesydx+Sgp/fjpuILIXlLJJ12X78J
1ikHXVk5efjG+ZMQ8pUYvIZHicuYw8mLJvUKpko6bZ3JnHI2PKJZnLG8tvv0n5HJyE9zVT06BxQw
ECDQBhYjibh+TuUjrRW7z3ye5bSYwOixyfeb4B5Fmb19oJsQg6ADwcgNhXxbzWWqgMffxyJVR7VI
QqRiye0e2XCPz7TAOlFXsYfKHIZ4xs4auhZLV+coT2sc/1WEv3Re1W/igp0QkeUepKn+NqCrHKHS
MBKdYFVbMpvc016FU9Vd+hDdwI6R/wX0D9sCJvpsAW24qv6861ZTPyo/s+5UVS9Mr3D9hlEflpsJ
NAJf3nDiJ/OwWgqa5eb+Jup1GX8Rmj+6fT/erduzIjU3yfcKpQv8vgB+a4DINZ9dovnV5RLdxq7q
muPt18TUrB+TnWHdtKq5A9St1j9pTiZ/or4vPuZWs2tr1cZzJm2qT/WiKlQaVYUz73p8uLdG53su
rhtphzvbGjTmKzf6/2rLYkuJUBWEFGx5oG9jML+IthYi5QHrLa4lP3YIHr8rXpNsx1b8vca3UT7X
3f22eWwGZnaqgkc29kND57fPyBN6wxj28CRKB12wJ2X/PH2CfNKy6GLEc2a+YXwt4EmPZXPk3Bge
d/lQ1864gvft21Pj84eaEMpXgq5F8G01pdWU45ZozbzFBoGg09bi5+r0R8hP51agFLiwPCrciOP8
J/8ZE/CrZmSc0DftutgIiPoBZEXd6ZXamKuuEu6kUbl1T8BcRVtXWlY+3zxKTgGNn1UC8ULElfD9
dMZLYcJZeYstxsq48rZsgXlAXBZmAfqbSjwL72OFz4b53y1YZCEZl63yASRdrGqt6TGHHJga6bqn
/XPNeSGtmbf8gRo20tP4IUw6psTKtgYRL1/hxrZ+xIHzij8CZzaXWhcA9d2LlyLjM2zywIt9Gd+U
6inpmhWmR7QBNj0ZtNqso7ilkkpUAmOVXwcowvRVO8ejid8rGLvOGIl0uw4EJ89yfgTyaJrj1OGS
Zk3iJa5HrI+s8nKYIWPf2yG5UV+IzaayR2kJ2A5zImdolQuCcUaYb/3QhbN/KSCrmb8ygHTompPd
KwdQtnp5nl4E6rWCPFfNb0eEJ3qkLm78uO30cmpK5qc4VTCc+4GYsmQrFonYEy+Zkm9zV+EGZtMG
46E1wrlmbj0kfNErCx8VhjTjqVQ5KRFpKU9MNG3CTnszmy/8zxnwumrEN0tsCQdhoIEBo7lSyV4C
/4rN5TafRocz1Dh9NP4JwcNO7bJLsRpEWauYyxMtq56oobkcWTZ+3MspiqmAmAEoWKcldkJlNgni
oFxvnEt4AH8rtwLvKnMWfe+lEHianTrVAIibNqRT5JX1XHelsqRTNVWxtvhXARkbOgUr6L1tbNdH
mhOOudhcSmcM5i0OxVX47irQzq+GvyXmzve8s2RVf4LPE3JjviFabzigNYFQcifGt0rQ53EBUyP+
Wusn1SMWKvlRjCXERUJByhMpklsNZXZ4r3SPj8lWVtkGHFbefseayqHTErQsDLh2iLDdRKiej0C9
oUnEq8zMf0sA3FelztREPZ/iixILuseUhkzsf9v+fA3WBflybtWbq5N9yiBF/yGcp6AOc39F86Lt
rs361IP4v7DGwlhcrfvF0ZkPwq69Bj18XVzMMX4mF4wm/RV+fJy8KLpRzE+5JaECpi6v7NuX3nom
4EaP/kRSIPzv53QQQcuaXW7d+xUfyZrdT+/EE5vRybB8ZfsGP+J/3tk4sfRc/zbXpcSORKMQvq22
nAm/KA7L5WVgNtPuDtKHkyvQHPnrOFeQ2uQZZQAyp3yNjNIK00Z1/jAhntaY/+rrcYLsqatQgixv
vtxyqbq1BhyugkPmRdWbvst9xJ9w1fQ6ByN5ZwzTfopmPF6oFfeMj+PD3j7Z6y7sT45fKhX7JDYt
VbrBSzXMpRrUm+pxIZMR0t1LWANQkwr5FLUj0F8PRXAhm/o1RAsdwQ5/YOh73nr1fvX9VmRRCkuw
GIqjtzRhykp24DD+pPbjjyOIa7o85irc3PtLJ7T3WKXFfYn4zpkAn+qIcjeGZeyieGFmMzlfQb3F
Y4CE4dX+DHB9obebHiX+z7p2VwD2N+joFSmlk6JEXfjA6NOIAPNIizlzmI605N6YldiEgxDP2Rnw
kLzdnSumy0bnogBgNfS4WKm53E/vNqkeS1XfvB8od7Jt/ZaSKgipR9+0LbZxf5lPJpYdqAJmf8In
W/kvGKfCadxAoci1As7A0iFEDVMqaGbMsdAud894bwjhe1T4ymjKeZym/QupMiNAyC7D3My/V/k5
2eVPDhe3e0F2Esei/2QF9GLRMh0pXuS2sKQQCN3YMvdc19FCZyX/S2yrhyTNP5Pcy+eGpXrE1EqC
jkvLO64hCiYSYOpNnpE0mu2NLoSvR9MpLM7QMGqMSbWJq/3fe9IubwPLIJGFeK0a1EX4HT/SQi39
kg14hQMYFy8zO+AAtB6/f71Kuo8cwUowA6cUCZxh+w31nwngtqJdrF5NnWBj0rTg6Kp1SAkYYuuB
5A9+wM3d9mYHEG3Z3InqaXIy0m35RLQxQr7JfxmwIr5lh/NdCjZOESSDZTvFgQuZG5JoCYGk1plk
gWcYVxGGM96PnmxVSF0ei0eKcG0KtfoWZ4eMtyTDEvkvzZhxWPOsGzFiLVNw71TMKbg33C05zC3D
Ot8ygcOjX9vBPaVka3ACSjxvF7KnQmCaW/ZfdE745EaSdk34kp8Rap2May30ouZJX12m7BGcdEIW
H7TVsBjsy2kr32ds3npg4hPtTsljlqe6PcFNpvm9HxCNf7o6YJ0YtroEJW2/r8BiWz3VmaHe9sJQ
0rcaGwTdehWyk9UbKJJyzQIX5A0RuYJWWbThWUKoj2dwU8jUF2TDViDz/yunEPBxm8w6I53eMQ2j
ccNtoOC6+JXKhId9XA7+nTuFP1bj+ipd+wisjCC7r7tKKRJjMzQEkO/BFfSAtJxS33xo+bK4t0K0
7X5k1q/RXH5O39woqoauVaOoXxmHc/4lfxlYkuaFj6P6PYGL6eqQBOsV18TFPioND4lFaMsUabmQ
hFVam4EDIbmLKRTtUCYX2Pp8YmLkqHsKrBqLjzPN7TGReCDvMmcV05PEXvjzBCxDcnOBoyyR7qUn
67MNJq5ePYuJ5d9k8+Zx5awUf75eOTwJm58PiPGN9zL8HxFSXtB1AulIAxQoxaC3gapXuLUSEMrM
++IvQVUczLGxsCrMprJqeON/ijEaZ9cIBGThF8g0WVGKSoQk/NsCBDk7UIXtPH0TEzUCgEAKbXp7
cVUzwVC7gP9GAwt/UH5NmpWYXrTyIjL+Nd+pQoq+rxPqflxP6/jLFjdtCPv3G5Koh7FRShEwJO0J
UrAFnVEJotXl4hv6MuXQfc7P1rjEOH110a3SaiyRKY1hd+FS+dw8dnYltT+pz3sEIJC0JBO5cXkK
CEdTkwwK7QvKE9w+R2WWpgU3gQZpzYoLdwz5VttEK4TAynxmSq6N2kuEKpK7R2TREbmEcpQTiRzn
IC0wFjcvpnwFU3D56VLrj+DqoRO7lY7UsIIxgXLhvfcTYivQmAkDGvGwpOr1SJ0QV7orP1xmeEt0
xvnZbHl6jrpF93wvcBtjw20zxNaChVNKSPY4PWe4i5mlGgm3MDZRickrzCUJN35WOURZ5OKU+5Px
nlWmKFvH07O3CbSb6dNdHAb/kZXez59hmyAJphStgjGRYv2TSFDEfCzS54uwHWW1n3RO1ClHAIk2
PVfRZsh6zWYmJNETE5CYnSimC9OQmUn50Z4brcohWfy4Z6tX2btSmN+WEgfiVo5FgftR4juqbdtt
EMHCZ7SCdwERohYJEkK/YIBYK2DDQBGL7bG1kRwlY5UFo0bKAO1DLE7pvRn34Ho1O7BzZgRk7V03
rI8+6GCrnueGevlAiehiOGHCpN4yhsK6zVPAZB3TAbSCMCv0IRAKk/vu8slQ9ZzIb7gDhz84QVjM
IHCJUuNU17z5+YW4biYaY+zfxdsOVfK7m0OZvNmpQG2Bs9zLOeSNz20zMysJ3o7JFUTXmFYlZJyO
aTVQ2BMOVXaHPEnQ03xos3fuSfPu291w76FHU71HV8HGnzJB7ZNVnyHUC5ppYa5Nwt3i+jJshw9P
RpYN3+ttXjw5U/R45ZMWVV/3AlUb2oaiSTWLVbQSzkbnAWAXrJ94mtDZnf/bU+h5MId1jajoC0U7
AZ/JwlXzYYcsnGtQaEUqiNApUkg+jOP8XaHWNQL3+wiAhBI3OrzqanACjO2GIBF9WtjaxraP8Gnb
rAZnUKZCt9RL+3PeO5xuDOX7ysaf5xAVjN4aHefcGgzEBW+//y677ZlS8b78UDdyvM21ijPmV0lv
Ae+FbsHfF4CO/Xn7o8CrqwtlYxBdgCve2/IpEYyOLeQYq1P/rRqshRwZBDip7mCYIjaKE0GbSeYH
057HMqlL7m3/1KBdEg3ajTkDJ5BiUMjwfveLBaTmHuQWY6h/EGFxbx9GIBxERE9jVkh0DlCnZGuh
wzTCf8Pkwfzq5YGQpykzntlgqrLvmRnRawMf2yExuIcHc1ljx6q5BB2bkm1mA31rvA1GfFIJtUNO
MbsOwj6SKKeUA+mM2pF2jlpSiWWZ9qw7lGWX5FSkZDgtOodmTPnxM6NC/E2TqEEweaLC8giQAAiW
ctfTuN1DKKqvt6n7ysxr5NgHUtBUnUJXaslftDFD/ri5S8MmQ763lP7mYCGpbJuSkJ9WOSqRa95A
Z+DGbMXx92N+vEWbOkPu9s/K/YOxnnpObfM99iDDuWDUMDgHr+pa+z7Jjy7nhuOW0C4tUjdy5kdn
YftjfgSuhh+2ZbYEEtx42moUJLe3yiWXEjadsjD/G1LNZn37ybkNNwOhCSCH0bD74EEhZRiSdusS
RkY1kEXFYKNuPBn3FuH8S0+hsJYlSk4Szo4/3m9zlWGdtJWlKyiA8yo0MJdzi9gomIdkveXkngpt
EL6b7SkbmLWWez2NLiwSda4Zbu94hlq9n8IuM4+StuQX2zPdSsQOb2y8SOcKT0VbzvlfW2r+j9uS
M3sj61Jpb0eyfX/UJDiCfK24NVRRxJHVc5CJBwac1yHX4WoFPqbtn+5P3z+SUCrB03YwSYluzf3H
MlZ6NmM2OtLnQX/KYSc8nTu6kY5Qyqd/dncmmxYfIC6Ub2pWmlPSDfyv+JdszyyI46AV8sbIrQhH
q2NXdT7TZYd8DN5wfY4ipsXWjiFJP+Ow4ThFlEfha3urX4494zEJH0EbB+de79frutvQIPphtdoQ
AyBUw/n/fPyMy3FMPPdTYRIBNfzYglIytyeLWBYcuXAuD6xlX83uyY+IyCdetTORl41wufIBUiP7
nWJDjJHl7HNFXnspaRA5U4/bPoVy80JdWOzOJgFaWXieJc2NS+ZlN+xt5461rnWqkE6gUGDS2ecK
fd57wBYnt73jSrFTfCvB0a6yIvAzvgTG0ec/tQ3ihlbx8GC+mnb3JUAR63ohuvG/JuMuDjU4CZWn
gLyX9jfZYjtTIg3MQcmsSCTMLK9qupzsveI7m7oSyW8nBf+zQKbi4Xms7YcwdES7DCTO1fNIAOtv
2+rmw+N5601bIBolXyYdjd5lUiUzDhmAOJCIG/BIqjzTjk6YXuxeV5563JCL8eLy/+hY4CuaWMxd
GSjn3Z/vdspSWDwcoMUsV2ivNL/5Ta/pTx3Jd+2gCn7E99EuuyhlzMSbtLifiDkNi9bPvJMW0mAB
TTmRlF6npEMCOtaMEz4P1YPorwVpTH+jFZTHYlrsn0ZTYHDI2lOT39f7Bcvvb0UflUF6TCGBHisv
rhC/FGwjJEezzvRvYsfeyONAWxO7Zy6gMoBrHll1/eB0KNA/DOTZmsQ6Ugj6SeqXU80Bw5rGxNkU
TlDBxtnMQT97YkTZycPjom9wg8p3EzTC8Xz8cR8WWWmlNLHFCLz6DTm+nTdLYReyKk5tAJZqo2F5
n7D+juG0drDbfkXyA3rTwA8me4hQ8rz9PbFqSIMjXOL1clsD3Q3ucJZ9Mt9gUJ0iaBMHaontGe5x
zUC085IvEduLzp1jes2hh2RZtRvrt36t/AywrqB9sEUN4W2mk2s/BD3JcjPQ8j90p2FLrBqEntoP
ymKo/hARZBG5EAZq1gQz51D5Y5PWNH12t+OhLe84gxFASJhpgVEZcZJ64BlnFODzuIKOj+FBD45c
KJVMMQTsmpYZ+IO4EvfFx5vjJ5g=
`pragma protect end_protected
module usb_fifo (
  Data,
  WrClk,
  RdClk,
  WrEn,
  RdEn,
  Almost_Empty,
  Almost_Full,
  Q,
  Empty,
  Full
)
;
input [7:0] Data;
input WrClk;
input RdClk;
input WrEn;
input RdEn;
output Almost_Empty;
output Almost_Full;
output [7:0] Q;
output Empty;
output Full;
wire VCC;
wire GND;
  \~fifo.usb_fifo  fifo_inst (
    .RdClk(RdClk),
    .WrClk(WrClk),
    .WrEn(WrEn),
    .RdEn(RdEn),
    .Data(Data[7:0]),
    .Full(Full),
    .Almost_Empty(Almost_Empty),
    .Almost_Full(Almost_Full),
    .Empty(Empty),
    .Q(Q[7:0])
);
  VCC VCC_cZ (
    .V(VCC)
);
  GND GND_cZ (
    .G(GND)
);
  GSR GSR (
    .GSRI(VCC) 
);
endmodule /* usb_fifo */

module ACMRequestHandlers(request, data_requested, status_requested, rx_ready_for_response, valid, ack, stall, last, \type );
  reg \$auto$verilog_backend.cc:2083:dump_module$1  = 0;
  wire \$1 ;
  wire \$3 ;
  wire \$5 ;
  wire \$7 ;
  wire \$9 ;
  output ack;
  reg ack;
  input data_requested;
  wire data_requested;
  output last;
  reg last;
  input [7:0] request;
  wire [7:0] request;
  input rx_ready_for_response;
  wire rx_ready_for_response;
  output stall;
  reg stall;
  input status_requested;
  wire status_requested;
  input [1:0] \type ;
  wire [1:0] \type ;
  output valid;
  reg valid;
  assign \$9  = status_requested |  data_requested;
  assign \$1  = \type  ==  1'h1;
  assign \$3  = \type  ==  1'h1;
  assign \$5  = \type  ==  1'h1;
  assign \$7  = \type  ==  1'h1;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    ack = 1'h0;
    casez (\$1 )
      1'h1:
          casez (request)
            8'h20:
                casez (rx_ready_for_response)
                  1'h1:
                      ack = 1'h1;
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    valid = 1'h0;
    casez (\$3 )
      1'h1:
          casez (request)
            8'h20:
                casez (status_requested)
                  1'h1:
                      valid = 1'h1;
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    last = 1'h0;
    casez (\$5 )
      1'h1:
          casez (request)
            8'h20:
                casez (status_requested)
                  1'h1:
                      last = 1'h1;
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    stall = 1'h0;
    casez (\$7 )
      1'h1:
          casez (request)
            8'h20:
                ;
            default:
                casez (\$9 )
                  1'h1:
                      stall = 1'h1;
                endcase
          endcase
    endcase
  end
endmodule
module StallOnlyRequestHandler(data_requested, status_requested, stall, \type );
  reg \$auto$verilog_backend.cc:2083:dump_module$2  = 0;
  wire \$1 ;
  wire \$3 ;
  wire \$5 ;
  wire \$7 ;
  input data_requested;
  wire data_requested;
  output stall;
  reg stall;
  input status_requested;
  wire status_requested;
  input [1:0] \type ;
  wire [1:0] \type ;
  assign \$1  = data_requested |  status_requested;
  assign \$3  = \type  ==  2'h2;
  assign \$5  = \type  ==  2'h3;
  assign \$7  = \$3  |  \$5 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$2 ) begin end
    stall = 1'h0;
    casez (\$1 )
      1'h1:
          casez (\$7 )
            1'h1:
                stall = 1'h1;
          endcase
    endcase
  end
endmodule
module StandardRequestHandler(usb_clk, \type , request, value, length, received, data_requested, status_requested, ack, active_config, address_changed, new_address, config_changed, new_config, valid, tx_data_pid, \ack$1 , stall, payload, first, last
, ready, usb_rst);
  reg \$auto$verilog_backend.cc:2083:dump_module$3  = 0;
  wire \$11 ;
  wire \$13 ;
  wire \$15 ;
  wire \$17 ;
  wire \$19 ;
  wire \$2 ;
  wire \$21 ;
  wire \$23 ;
  wire \$25 ;
  wire \$27 ;
  wire \$29 ;
  wire \$31 ;
  wire \$33 ;
  wire \$35 ;
  wire \$37 ;
  wire \$39 ;
  wire \$4 ;
  wire \$41 ;
  wire \$43 ;
  wire \$45 ;
  wire \$47 ;
  wire \$49 ;
  wire [7:0] \$51 ;
  wire \$53 ;
  wire \$55 ;
  wire \$57 ;
  wire \$59 ;
  wire [11:0] \$6 ;
  wire [11:0] \$7 ;
  wire \$9 ;
  input ack;
  wire ack;
  output \ack$1 ;
  reg \ack$1 ;
  input [7:0] active_config;
  wire [7:0] active_config;
  output address_changed;
  reg address_changed;
  output config_changed;
  reg config_changed;
  input data_requested;
  wire data_requested;
  reg expecting_ack = 1'h0;
  reg \expecting_ack$next ;
  output first;
  reg first;
  reg [2:0] fsm_state = 3'h0;
  reg [2:0] \fsm_state$next ;
  wire get_descriptor_first;
  wire get_descriptor_last;
  wire [15:0] get_descriptor_length;
  wire [7:0] get_descriptor_payload;
  reg get_descriptor_ready;
  wire get_descriptor_stall;
  reg get_descriptor_start;
  reg [10:0] get_descriptor_start_position = 11'h000;
  reg [10:0] \get_descriptor_start_position$next ;
  wire get_descriptor_valid;
  wire [15:0] get_descriptor_value;
  output last;
  reg last;
  input [15:0] length;
  wire [15:0] length;
  output [6:0] new_address;
  reg [6:0] new_address;
  output [7:0] new_config;
  reg [7:0] new_config;
  output [7:0] payload;
  reg [7:0] payload;
  input ready;
  wire ready;
  input received;
  wire received;
  input [7:0] request;
  wire [7:0] request;
  output stall;
  reg stall;
  input status_requested;
  wire status_requested;
  reg [7:0] transmitter_datum_0;
  reg [7:0] transmitter_datum_1;
  wire transmitter_first;
  wire transmitter_last;
  reg [1:0] transmitter_max_length;
  wire [7:0] transmitter_payload;
  reg transmitter_ready;
  reg transmitter_start;
  wire transmitter_valid;
  output tx_data_pid;
  reg tx_data_pid = 1'h1;
  reg \tx_data_pid$next ;
  input [1:0] \type ;
  wire [1:0] \type ;
  input usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  output valid;
  reg valid;
  input [15:0] value;
  wire [15:0] value;
  assign \$9  = !  \type ;
  assign \$11  = ack &  expecting_ack;
  assign \$13  = ~  tx_data_pid;
  assign \$15  = !  \type ;
  assign \$19  = data_requested |  status_requested;
  assign \$21  = !  \type ;
  assign \$23  = !  \type ;
  assign \$25  = !  \type ;
  assign \$27  = !  \type ;
  assign \$2  = !  \type ;
  assign \$29  = !  \type ;
  assign \$31  = !  \type ;
  assign \$33  = !  \type ;
  assign \$35  = !  \type ;
  assign \$37  = !  \type ;
  assign \$39  = !  \type ;
  assign \$41  = data_requested |  status_requested;
  assign \$43  = !  \type ;
  assign \$45  = !  \type ;
  assign \$47  = !  \type ;
  assign \$4  = ack &  expecting_ack;
  assign \$49  = !  \type ;
  assign \$51  = +  value[6:0];
  assign \$53  = !  \type ;
  assign \$55  = !  \type ;
  assign \$57  = !  \type ;
  assign \$59  = ack &  expecting_ack;
  always @(posedge usb_clk)
    get_descriptor_start_position <= \get_descriptor_start_position$next ;
  always @(posedge usb_clk)
    tx_data_pid <= \tx_data_pid$next ;
  always @(posedge usb_clk)
    fsm_state <= \fsm_state$next ;
  always @(posedge usb_clk)
    expecting_ack <= \expecting_ack$next ;
  assign \$7  = get_descriptor_start_position +  7'h40;
  get_descriptor get_descriptor (
    .first(get_descriptor_first),
    .last(get_descriptor_last),
    .length(get_descriptor_length),
    .payload(get_descriptor_payload),
    .ready(get_descriptor_ready),
    .stall(get_descriptor_stall),
    .start(get_descriptor_start),
    .start_position(get_descriptor_start_position),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst),
    .valid(get_descriptor_valid),
    .value(get_descriptor_value)
  );
  \transmitter$4  transmitter (
    .datum_0(transmitter_datum_0),
    .datum_1(transmitter_datum_1),
    .first(transmitter_first),
    .last(transmitter_last),
    .max_length(transmitter_max_length),
    .payload(transmitter_payload),
    .ready(transmitter_ready),
    .start(transmitter_start),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst),
    .valid(transmitter_valid)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    transmitter_datum_0 = 8'h00;
    transmitter_datum_1 = 8'h00;
    casez (\$31 )
      1'h1:
          casez (fsm_state)
            3'h0:
                ;
            3'h1:
                { transmitter_datum_1, transmitter_datum_0 } = 16'h0000;
            3'h2:
                ;
            3'h3:
                ;
            3'h4:
                ;
            3'h5:
                transmitter_datum_0 = active_config;
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    transmitter_max_length = 2'h0;
    casez (\$33 )
      1'h1:
          casez (fsm_state)
            3'h0:
                ;
            3'h1:
                transmitter_max_length = 2'h2;
            3'h2:
                ;
            3'h3:
                ;
            3'h4:
                ;
            3'h5:
                transmitter_max_length = 2'h1;
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    transmitter_start = 1'h0;
    casez (\$35 )
      1'h1:
          casez (fsm_state)
            3'h0:
                ;
            3'h1:
                casez (data_requested)
                  1'h1:
                      transmitter_start = 1'h1;
                endcase
            3'h2:
                ;
            3'h3:
                ;
            3'h4:
                ;
            3'h5:
                casez (data_requested)
                  1'h1:
                      transmitter_start = 1'h1;
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    \ack$1  = 1'h0;
    casez (\$37 )
      1'h1:
          casez (fsm_state)
            3'h0:
                ;
            3'h1:
                casez (status_requested)
                  1'h1:
                      \ack$1  = 1'h1;
                endcase
            3'h2:
                ;
            3'h3:
                ;
            3'h4:
                casez (status_requested)
                  1'h1:
                      \ack$1  = 1'h1;
                endcase
            3'h5:
                casez (status_requested)
                  1'h1:
                      \ack$1  = 1'h1;
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    stall = 1'h0;
    casez (\$39 )
      1'h1:
          casez (fsm_state)
            3'h0:
                ;
            3'h1:
                ;
            3'h2:
                ;
            3'h3:
                ;
            3'h4:
                stall = get_descriptor_stall;
            3'h5:
                ;
            3'h6:
                casez (\$41 )
                  1'h1:
                      stall = 1'h1;
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    address_changed = 1'h0;
    casez (\$43 )
      1'h1:
          casez (fsm_state)
            3'h0:
                ;
            3'h1:
                ;
            3'h2:
                casez (ack)
                  1'h1:
                      address_changed = 1'h1;
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    new_address = 7'h00;
    casez (\$45 )
      1'h1:
          casez (fsm_state)
            3'h0:
                ;
            3'h1:
                ;
            3'h2:
                casez (ack)
                  1'h1:
                      new_address = value[6:0];
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    config_changed = 1'h0;
    casez (\$47 )
      1'h1:
          casez (fsm_state)
            3'h0:
                ;
            3'h1:
                ;
            3'h2:
                ;
            3'h3:
                casez (ack)
                  1'h1:
                      config_changed = 1'h1;
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    new_config = 8'h00;
    casez (\$49 )
      1'h1:
          casez (fsm_state)
            3'h0:
                ;
            3'h1:
                ;
            3'h2:
                ;
            3'h3:
                casez (ack)
                  1'h1:
                      new_config = \$51 ;
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    \get_descriptor_start_position$next  = get_descriptor_start_position;
    casez (\$2 )
      1'h1:
          casez (fsm_state)
            3'h0:
                \get_descriptor_start_position$next  = 11'h000;
            3'h1:
                ;
            3'h2:
                ;
            3'h3:
                ;
            3'h4:
                casez (\$4 )
                  1'h1:
                      \get_descriptor_start_position$next  = \$7 [10:0];
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \get_descriptor_start_position$next  = 11'h000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    get_descriptor_ready = 1'h0;
    casez (\$53 )
      1'h1:
          casez (fsm_state)
            3'h0:
                ;
            3'h1:
                ;
            3'h2:
                ;
            3'h3:
                ;
            3'h4:
                get_descriptor_ready = ready;
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    get_descriptor_start = 1'h0;
    casez (\$55 )
      1'h1:
          casez (fsm_state)
            3'h0:
                ;
            3'h1:
                ;
            3'h2:
                ;
            3'h3:
                ;
            3'h4:
                casez (data_requested)
                  1'h1:
                      get_descriptor_start = 1'h1;
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    \expecting_ack$next  = expecting_ack;
    casez (\$57 )
      1'h1:
          casez (fsm_state)
            3'h0:
                ;
            3'h1:
                ;
            3'h2:
                ;
            3'h3:
                ;
            3'h4:
              begin
                casez (data_requested)
                  1'h1:
                      \expecting_ack$next  = 1'h1;
                endcase
                casez (\$59 )
                  1'h1:
                      \expecting_ack$next  = 1'h0;
                endcase
              end
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \expecting_ack$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    \tx_data_pid$next  = tx_data_pid;
    casez (\$9 )
      1'h1:
          casez (fsm_state)
            3'h0:
                \tx_data_pid$next  = 1'h1;
            3'h1:
                ;
            3'h2:
                ;
            3'h3:
                ;
            3'h4:
                casez (\$11 )
                  1'h1:
                      \tx_data_pid$next  = \$13 ;
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \tx_data_pid$next  = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    \fsm_state$next  = fsm_state;
    casez (\$15 )
      1'h1:
          casez (fsm_state)
            3'h0:
                casez (received)
                  1'h1:
                      casez (\$17 )
                        1'h1:
                            casez (request)
                              8'h00:
                                  \fsm_state$next  = 3'h1;
                              8'h05:
                                  \fsm_state$next  = 3'h2;
                              8'h09:
                                  \fsm_state$next  = 3'h3;
                              8'h06:
                                  \fsm_state$next  = 3'h4;
                              8'h08:
                                  \fsm_state$next  = 3'h5;
                              default:
                                  \fsm_state$next  = 3'h6;
                            endcase
                      endcase
                endcase
            3'h1:
                casez (status_requested)
                  1'h1:
                      \fsm_state$next  = 3'h0;
                endcase
            3'h2:
                casez (ack)
                  1'h1:
                      \fsm_state$next  = 3'h0;
                endcase
            3'h3:
                casez (ack)
                  1'h1:
                      \fsm_state$next  = 3'h0;
                endcase
            3'h4:
                casez (status_requested)
                  1'h1:
                      \fsm_state$next  = 3'h0;
                endcase
            3'h5:
                casez (status_requested)
                  1'h1:
                      \fsm_state$next  = 3'h0;
                endcase
            3'h6:
                casez (\$19 )
                  1'h1:
                      \fsm_state$next  = 3'h0;
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \fsm_state$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    valid = 1'h0;
    casez (\$21 )
      1'h1:
          casez (fsm_state)
            3'h0:
                ;
            3'h1:
                valid = transmitter_valid;
            3'h2:
                casez (status_requested)
                  1'h1:
                      valid = 1'h1;
                endcase
            3'h3:
                casez (status_requested)
                  1'h1:
                      valid = 1'h1;
                endcase
            3'h4:
                valid = get_descriptor_valid;
            3'h5:
                valid = transmitter_valid;
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    first = 1'h0;
    casez (\$23 )
      1'h1:
          casez (fsm_state)
            3'h0:
                ;
            3'h1:
                first = transmitter_first;
            3'h2:
                ;
            3'h3:
                ;
            3'h4:
                first = get_descriptor_first;
            3'h5:
                first = transmitter_first;
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    last = 1'h0;
    casez (\$25 )
      1'h1:
          casez (fsm_state)
            3'h0:
                ;
            3'h1:
                last = transmitter_last;
            3'h2:
                casez (status_requested)
                  1'h1:
                      last = 1'h1;
                endcase
            3'h3:
                casez (status_requested)
                  1'h1:
                      last = 1'h1;
                endcase
            3'h4:
                last = get_descriptor_last;
            3'h5:
                last = transmitter_last;
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    payload = 8'h00;
    casez (\$27 )
      1'h1:
          casez (fsm_state)
            3'h0:
                ;
            3'h1:
                payload = transmitter_payload;
            3'h2:
                ;
            3'h3:
                ;
            3'h4:
                payload = get_descriptor_payload;
            3'h5:
                payload = transmitter_payload;
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    transmitter_ready = 1'h0;
    casez (\$29 )
      1'h1:
          casez (fsm_state)
            3'h0:
                ;
            3'h1:
                transmitter_ready = ready;
            3'h2:
                ;
            3'h3:
                ;
            3'h4:
                ;
            3'h5:
                transmitter_ready = ready;
          endcase
    endcase
  end
  assign \$6  = \$7 ;
  assign get_descriptor_length = length;
  assign get_descriptor_value = value;
  assign \$17  = 1'h1;
endmodule
module USBControlEndpoint(rx_valid, usb_rst, usb_clk, rx_active, crc, tx_allowed, tx_timeout, rx_timeout, ack, nak, stall, nyet, pid, address, endpoint, new_token, ready_for_response, frame, new_frame, is_in, is_out
, is_setup, is_ping, valid, next, payload, rx_ready_for_response, speed, active_config, address_changed, new_address, config_changed, new_config, \ack$1 , \nak$2 , \stall$3 , start, \start$4 , \valid$5 , tx_pid_toggle, \payload$6 , first
, last, ready, rx_data);
  reg \$auto$verilog_backend.cc:2083:dump_module$4  = 0;
  wire \$100 ;
  wire \$102 ;
  wire \$104 ;
  wire \$106 ;
  wire \$108 ;
  wire \$110 ;
  wire \$112 ;
  wire \$114 ;
  wire \$116 ;
  wire \$118 ;
  wire \$120 ;
  wire \$122 ;
  wire \$124 ;
  wire \$126 ;
  wire \$128 ;
  wire \$130 ;
  wire \$132 ;
  wire \$134 ;
  wire \$58 ;
  wire \$60 ;
  wire \$62 ;
  wire \$64 ;
  wire \$66 ;
  wire \$68 ;
  wire \$70 ;
  wire [1:0] \$72 ;
  wire \$74 ;
  wire \$76 ;
  wire \$78 ;
  wire \$80 ;
  wire \$82 ;
  wire \$84 ;
  wire \$86 ;
  wire \$88 ;
  wire \$90 ;
  wire \$92 ;
  wire \$94 ;
  wire \$96 ;
  wire \$98 ;
  input ack;
  wire ack;
  output \ack$1 ;
  reg \ack$1 ;
  input [7:0] active_config;
  wire [7:0] active_config;
  input [6:0] address;
  wire [6:0] address;
  wire [6:0] \address$47 ;
  output address_changed;
  wire address_changed;
  output config_changed;
  wire config_changed;
  input [15:0] crc;
  wire [15:0] crc;
  input [3:0] endpoint;
  wire [3:0] endpoint;
  wire [3:0] \endpoint$48 ;
  output first;
  wire first;
  input [10:0] frame;
  wire [10:0] frame;
  wire [10:0] \frame$50 ;
  reg [2:0] fsm_state = 3'h0;
  reg [2:0] \fsm_state$next ;
  input is_in;
  wire is_in;
  wire \is_in$52 ;
  input is_out;
  wire is_out;
  wire \is_out$53 ;
  input is_ping;
  wire is_ping;
  wire \is_ping$55 ;
  input is_setup;
  wire is_setup;
  wire \is_setup$54 ;
  output last;
  wire last;
  input nak;
  wire nak;
  output \nak$2 ;
  wire \nak$2 ;
  output [6:0] new_address;
  wire [6:0] new_address;
  output [7:0] new_config;
  wire [7:0] new_config;
  input new_frame;
  wire new_frame;
  wire \new_frame$51 ;
  input new_token;
  wire new_token;
  input next;
  wire next;
  input nyet;
  wire nyet;
  input [7:0] payload;
  wire [7:0] payload;
  output [7:0] \payload$6 ;
  wire [7:0] \payload$6 ;
  input [3:0] pid;
  wire [3:0] pid;
  input ready;
  wire ready;
  input ready_for_response;
  wire ready_for_response;
  wire \ready_for_response$49 ;
  wire request_mux_ack;
  wire \request_mux_ack$20 ;
  wire \request_mux_ack$37 ;
  wire \request_mux_ack$38 ;
  wire \request_mux_ack$8 ;
  wire [7:0] request_mux_active_config;
  wire [7:0] \request_mux_active_config$21 ;
  wire [6:0] request_mux_address;
  wire request_mux_address_changed;
  wire \request_mux_address_changed$30 ;
  wire request_mux_config_changed;
  wire \request_mux_config_changed$32 ;
  reg request_mux_data_requested;
  wire \request_mux_data_requested$18 ;
  wire \request_mux_data_requested$24 ;
  wire \request_mux_data_requested$28 ;
  wire [3:0] request_mux_endpoint;
  wire request_mux_first;
  wire \request_mux_first$43 ;
  wire [10:0] request_mux_frame;
  wire [15:0] request_mux_index;
  wire request_mux_is_in;
  wire request_mux_is_in_request;
  wire request_mux_is_out;
  wire request_mux_is_ping;
  wire request_mux_is_setup;
  wire request_mux_last;
  wire \request_mux_last$44 ;
  wire \request_mux_last$45 ;
  wire [15:0] request_mux_length;
  wire [15:0] \request_mux_length$16 ;
  wire request_mux_nak;
  wire \request_mux_nak$9 ;
  wire [6:0] request_mux_new_address;
  wire [6:0] \request_mux_new_address$31 ;
  wire [7:0] request_mux_new_config;
  wire [7:0] \request_mux_new_config$33 ;
  wire request_mux_new_frame;
  wire request_mux_new_token;
  reg request_mux_next;
  wire request_mux_nyet;
  wire [7:0] request_mux_payload;
  reg [7:0] \request_mux_payload$12 ;
  wire [7:0] \request_mux_payload$42 ;
  wire [3:0] request_mux_pid;
  wire request_mux_ready;
  wire \request_mux_ready$46 ;
  wire request_mux_ready_for_response;
  wire request_mux_received;
  wire \request_mux_received$17 ;
  wire [4:0] request_mux_recipient;
  wire [7:0] request_mux_request;
  wire [7:0] \request_mux_request$14 ;
  wire [7:0] \request_mux_request$23 ;
  reg request_mux_rx_ready_for_response;
  wire \request_mux_rx_ready_for_response$26 ;
  wire request_mux_stall;
  wire \request_mux_stall$10 ;
  wire \request_mux_stall$39 ;
  wire \request_mux_stall$40 ;
  wire \request_mux_stall$41 ;
  reg request_mux_status_requested;
  wire \request_mux_status_requested$19 ;
  wire \request_mux_status_requested$25 ;
  wire \request_mux_status_requested$29 ;
  wire request_mux_tx_data_pid;
  wire \request_mux_tx_data_pid$35 ;
  wire [1:0] request_mux_type;
  wire [1:0] \request_mux_type$13 ;
  wire [1:0] \request_mux_type$22 ;
  wire [1:0] \request_mux_type$27 ;
  wire request_mux_valid;
  reg \request_mux_valid$11 ;
  wire \request_mux_valid$34 ;
  wire \request_mux_valid$36 ;
  wire [15:0] request_mux_value;
  wire [15:0] \request_mux_value$15 ;
  input rx_active;
  wire rx_active;
  input [7:0] rx_data;
  wire [7:0] rx_data;
  input rx_ready_for_response;
  wire rx_ready_for_response;
  input rx_timeout;
  wire rx_timeout;
  wire \rx_timeout$57 ;
  input rx_valid;
  wire rx_valid;
  wire setup_decoder_ack;
  wire [15:0] setup_decoder_crc;
  wire [15:0] setup_decoder_index;
  wire setup_decoder_is_in_request;
  wire [15:0] setup_decoder_length;
  wire setup_decoder_new_token;
  wire [3:0] setup_decoder_pid;
  wire setup_decoder_received;
  wire [4:0] setup_decoder_recipient;
  wire [7:0] setup_decoder_request;
  wire [1:0] setup_decoder_speed;
  wire setup_decoder_start;
  wire \setup_decoder_start$7 ;
  wire setup_decoder_tx_allowed;
  wire [1:0] setup_decoder_type;
  wire [15:0] setup_decoder_value;
  input [1:0] speed;
  wire [1:0] speed;
  input stall;
  wire stall;
  output \stall$3 ;
  wire \stall$3 ;
  output start;
  wire start;
  output \start$4 ;
  wire \start$4 ;
  input tx_allowed;
  wire tx_allowed;
  output [1:0] tx_pid_toggle;
  wire [1:0] tx_pid_toggle;
  input tx_timeout;
  wire tx_timeout;
  wire \tx_timeout$56 ;
  input usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  input valid;
  wire valid;
  output \valid$5 ;
  wire \valid$5 ;
  assign \$100  = new_token &  is_setup;
  assign \$102  = !  endpoint;
  assign \$104  = ready_for_response &  \$102 ;
  assign \$106  = \$104  &  is_in;
  assign \$108  = !  endpoint;
  assign \$110  = \$108  &  is_out;
  assign \$112  = !  endpoint;
  assign \$114  = \$112  &  is_out;
  assign \$116  = !  endpoint;
  assign \$118  = \$116  &  is_out;
  assign \$120  = !  endpoint;
  assign \$122  = \$120  &  is_out;
  assign \$124  = !  endpoint;
  assign \$126  = ready_for_response &  \$124 ;
  assign \$128  = \$126  &  is_in;
  assign \$130  = !  endpoint;
  assign \$132  = rx_ready_for_response &  \$130 ;
  assign \$134  = \$132  &  is_out;
  always @(posedge usb_clk)
    fsm_state <= \fsm_state$next ;
  assign \$58  = setup_decoder_ack |  request_mux_ack;
  assign \$60  = !  endpoint;
  assign \$62  = \$60  &  ready_for_response;
  assign \$64  = \$62  &  is_ping;
  assign \$66  = !  endpoint;
  assign \$68  = \$66  &  ready_for_response;
  assign \$70  = \$68  &  is_ping;
  assign \$72  = +  request_mux_tx_data_pid;
  assign \$74  = !  endpoint;
  assign \$76  = setup_decoder_received &  \$74 ;
  assign \$78  = |  setup_decoder_length;
  assign \$80  = new_token &  is_setup;
  assign \$82  = !  endpoint;
  assign \$84  = \$82  &  new_token;
  assign \$86  = is_out |  is_ping;
  assign \$88  = \$84  &  \$86 ;
  assign \$90  = new_token &  is_setup;
  assign \$92  = !  endpoint;
  assign \$94  = \$92  &  new_token;
  assign \$96  = \$94  &  is_in;
  assign \$98  = new_token &  is_setup;
  ACMRequestHandlers ACMRequestHandlers (
    .ack(\request_mux_ack$38 ),
    .data_requested(\request_mux_data_requested$24 ),
    .last(\request_mux_last$45 ),
    .request(\request_mux_request$23 ),
    .rx_ready_for_response(\request_mux_rx_ready_for_response$26 ),
    .stall(\request_mux_stall$40 ),
    .status_requested(\request_mux_status_requested$25 ),
    .\type (\request_mux_type$22 ),
    .valid(\request_mux_valid$36 )
  );
  StallOnlyRequestHandler StallOnlyRequestHandler (
    .data_requested(\request_mux_data_requested$28 ),
    .stall(\request_mux_stall$41 ),
    .status_requested(\request_mux_status_requested$29 ),
    .\type (\request_mux_type$27 )
  );
  StandardRequestHandler StandardRequestHandler (
    .ack(\request_mux_ack$20 ),
    .\ack$1 (\request_mux_ack$37 ),
    .active_config(\request_mux_active_config$21 ),
    .address_changed(\request_mux_address_changed$30 ),
    .config_changed(\request_mux_config_changed$32 ),
    .data_requested(\request_mux_data_requested$18 ),
    .first(\request_mux_first$43 ),
    .last(\request_mux_last$44 ),
    .length(\request_mux_length$16 ),
    .new_address(\request_mux_new_address$31 ),
    .new_config(\request_mux_new_config$33 ),
    .payload(\request_mux_payload$42 ),
    .ready(\request_mux_ready$46 ),
    .received(\request_mux_received$17 ),
    .request(\request_mux_request$14 ),
    .stall(\request_mux_stall$39 ),
    .status_requested(\request_mux_status_requested$19 ),
    .tx_data_pid(\request_mux_tx_data_pid$35 ),
    .\type (\request_mux_type$13 ),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst),
    .valid(\request_mux_valid$34 ),
    .value(\request_mux_value$15 )
  );
  request_mux request_mux (
    .ack(request_mux_ack),
    .\ack$1 (\request_mux_ack$8 ),
    .\ack$13 (\request_mux_ack$20 ),
    .\ack$30 (\request_mux_ack$37 ),
    .\ack$31 (\request_mux_ack$38 ),
    .active_config(request_mux_active_config),
    .\active_config$14 (\request_mux_active_config$21 ),
    .address(request_mux_address),
    .address_changed(request_mux_address_changed),
    .\address_changed$23 (\request_mux_address_changed$30 ),
    .config_changed(request_mux_config_changed),
    .\config_changed$25 (\request_mux_config_changed$32 ),
    .data_requested(request_mux_data_requested),
    .\data_requested$11 (\request_mux_data_requested$18 ),
    .\data_requested$17 (\request_mux_data_requested$24 ),
    .\data_requested$21 (\request_mux_data_requested$28 ),
    .endpoint(request_mux_endpoint),
    .first(request_mux_first),
    .\first$36 (\request_mux_first$43 ),
    .frame(request_mux_frame),
    .index(request_mux_index),
    .is_in(request_mux_is_in),
    .is_in_request(request_mux_is_in_request),
    .is_out(request_mux_is_out),
    .is_ping(request_mux_is_ping),
    .is_setup(request_mux_is_setup),
    .last(request_mux_last),
    .\last$37 (\request_mux_last$44 ),
    .\last$38 (\request_mux_last$45 ),
    .length(request_mux_length),
    .\length$9 (\request_mux_length$16 ),
    .nak(request_mux_nak),
    .\nak$2 (\request_mux_nak$9 ),
    .new_address(request_mux_new_address),
    .\new_address$24 (\request_mux_new_address$31 ),
    .new_config(request_mux_new_config),
    .\new_config$26 (\request_mux_new_config$33 ),
    .new_frame(request_mux_new_frame),
    .new_token(request_mux_new_token),
    .next(request_mux_next),
    .nyet(request_mux_nyet),
    .payload(request_mux_payload),
    .\payload$35 (\request_mux_payload$42 ),
    .\payload$5 (\request_mux_payload$12 ),
    .pid(request_mux_pid),
    .ready(request_mux_ready),
    .\ready$39 (\request_mux_ready$46 ),
    .ready_for_response(request_mux_ready_for_response),
    .received(request_mux_received),
    .\received$10 (\request_mux_received$17 ),
    .recipient(request_mux_recipient),
    .request(request_mux_request),
    .\request$16 (\request_mux_request$23 ),
    .\request$7 (\request_mux_request$14 ),
    .rx_ready_for_response(request_mux_rx_ready_for_response),
    .\rx_ready_for_response$19 (\request_mux_rx_ready_for_response$26 ),
    .stall(request_mux_stall),
    .\stall$3 (\request_mux_stall$10 ),
    .\stall$32 (\request_mux_stall$39 ),
    .\stall$33 (\request_mux_stall$40 ),
    .\stall$34 (\request_mux_stall$41 ),
    .status_requested(request_mux_status_requested),
    .\status_requested$12 (\request_mux_status_requested$19 ),
    .\status_requested$18 (\request_mux_status_requested$25 ),
    .\status_requested$22 (\request_mux_status_requested$29 ),
    .tx_data_pid(request_mux_tx_data_pid),
    .\tx_data_pid$28 (\request_mux_tx_data_pid$35 ),
    .\type (request_mux_type),
    .\type$15 (\request_mux_type$22 ),
    .\type$20 (\request_mux_type$27 ),
    .\type$6 (\request_mux_type$13 ),
    .valid(request_mux_valid),
    .\valid$27 (\request_mux_valid$34 ),
    .\valid$29 (\request_mux_valid$36 ),
    .\valid$4 (\request_mux_valid$11 ),
    .value(request_mux_value),
    .\value$8 (\request_mux_value$15 )
  );
  setup_decoder setup_decoder (
    .ack(setup_decoder_ack),
    .crc(setup_decoder_crc),
    .index(setup_decoder_index),
    .is_in_request(setup_decoder_is_in_request),
    .length(setup_decoder_length),
    .new_token(setup_decoder_new_token),
    .pid(setup_decoder_pid),
    .received(setup_decoder_received),
    .recipient(setup_decoder_recipient),
    .request(setup_decoder_request),
    .rx_active(rx_active),
    .rx_data(rx_data),
    .rx_valid(rx_valid),
    .speed(setup_decoder_speed),
    .start(setup_decoder_start),
    .\start$1 (\setup_decoder_start$7 ),
    .tx_allowed(setup_decoder_tx_allowed),
    .\type (setup_decoder_type),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst),
    .value(setup_decoder_value)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$4 ) begin end
    \ack$1  = \$58 ;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          casez (\$64 )
            1'h1:
                \ack$1  = 1'h1;
          endcase
      3'h3:
          ;
      3'h4:
          casez (\$70 )
            1'h1:
                \ack$1  = 1'h1;
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$4 ) begin end
    \fsm_state$next  = fsm_state;
    casez (fsm_state)
      3'h0:
          casez (\$76 )
            1'h1:
                casez (\$78 )
                  1'h1:
                      casez (setup_decoder_is_in_request)
                        1'h1:
                            \fsm_state$next  = 3'h1;
                        default:
                            \fsm_state$next  = 3'h2;
                      endcase
                  default:
                      \fsm_state$next  = 3'h3;
                endcase
          endcase
      3'h1:
        begin
          casez (\$80 )
            1'h1:
                \fsm_state$next  = 3'h0;
          endcase
          casez (\$88 )
            1'h1:
                \fsm_state$next  = 3'h4;
          endcase
        end
      3'h2:
        begin
          casez (\$90 )
            1'h1:
                \fsm_state$next  = 3'h0;
          endcase
          casez (\$96 )
            1'h1:
                \fsm_state$next  = 3'h3;
          endcase
        end
      3'h3:
          casez (\$98 )
            1'h1:
                \fsm_state$next  = 3'h0;
          endcase
      3'h4:
          casez (\$100 )
            1'h1:
                \fsm_state$next  = 3'h0;
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \fsm_state$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$4 ) begin end
    request_mux_data_requested = 1'h0;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          casez (\$106 )
            1'h1:
                request_mux_data_requested = 1'h1;
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$4 ) begin end
    \request_mux_valid$11  = 1'h0;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          casez (\$110 )
            1'h1:
                \request_mux_valid$11  = valid;
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$4 ) begin end
    request_mux_next = 1'h0;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          casez (\$114 )
            1'h1:
                request_mux_next = next;
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$4 ) begin end
    \request_mux_payload$12  = 8'h00;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          casez (\$118 )
            1'h1:
                \request_mux_payload$12  = payload;
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$4 ) begin end
    request_mux_rx_ready_for_response = 1'h0;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          casez (\$122 )
            1'h1:
                request_mux_rx_ready_for_response = rx_ready_for_response;
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$4 ) begin end
    request_mux_status_requested = 1'h0;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          ;
      3'h3:
          casez (\$128 )
            1'h1:
                request_mux_status_requested = 1'h1;
          endcase
      3'h4:
          casez (\$134 )
            1'h1:
                request_mux_status_requested = 1'h1;
          endcase
    endcase
  end
  assign tx_pid_toggle = \$72 ;
  assign new_config = request_mux_new_config;
  assign config_changed = request_mux_config_changed;
  assign request_mux_active_config = active_config;
  assign new_address = request_mux_new_address;
  assign address_changed = request_mux_address_changed;
  assign request_mux_nyet = nyet;
  assign \request_mux_stall$10  = stall;
  assign \request_mux_nak$9  = nak;
  assign \request_mux_ack$8  = ack;
  assign \stall$3  = request_mux_stall;
  assign \nak$2  = request_mux_nak;
  assign request_mux_ready = ready;
  assign \payload$6  = request_mux_payload;
  assign last = request_mux_last;
  assign first = request_mux_first;
  assign \valid$5  = request_mux_valid;
  assign request_mux_is_ping = is_ping;
  assign request_mux_is_setup = is_setup;
  assign request_mux_is_out = is_out;
  assign request_mux_is_in = is_in;
  assign request_mux_new_frame = new_frame;
  assign request_mux_frame = frame;
  assign request_mux_ready_for_response = ready_for_response;
  assign request_mux_new_token = new_token;
  assign request_mux_endpoint = endpoint;
  assign request_mux_address = address;
  assign request_mux_pid = pid;
  assign request_mux_received = setup_decoder_received;
  assign request_mux_length = setup_decoder_length;
  assign request_mux_index = setup_decoder_index;
  assign request_mux_value = setup_decoder_value;
  assign request_mux_request = setup_decoder_request;
  assign request_mux_is_in_request = setup_decoder_is_in_request;
  assign request_mux_type = setup_decoder_type;
  assign request_mux_recipient = setup_decoder_recipient;
  assign \start$4  = \setup_decoder_start$7 ;
  assign \rx_timeout$57  = rx_timeout;
  assign \tx_timeout$56  = tx_timeout;
  assign setup_decoder_tx_allowed = tx_allowed;
  assign setup_decoder_speed = speed;
  assign \is_ping$55  = is_ping;
  assign \is_setup$54  = is_setup;
  assign \is_out$53  = is_out;
  assign \is_in$52  = is_in;
  assign \new_frame$51  = new_frame;
  assign \frame$50  = frame;
  assign \ready_for_response$49  = ready_for_response;
  assign setup_decoder_new_token = new_token;
  assign \endpoint$48  = endpoint;
  assign \address$47  = address;
  assign setup_decoder_pid = pid;
  assign setup_decoder_crc = crc;
  assign start = setup_decoder_start;
endmodule
module USBStreamInEndpoint(usb_clk, ack, nak, stall, nyet, pid, address, endpoint, new_token, ready_for_response, frame, new_frame, is_in, is_out, is_setup, is_ping, \ack$1 , \nak$2 , \stall$3 , valid, tx_pid_toggle
, payload, first, last, ready, usb_rst);
  wire \$8 ;
  input ack;
  wire ack;
  output \ack$1 ;
  wire \ack$1 ;
  wire \ack$24 ;
  input [6:0] address;
  wire [6:0] address;
  wire [6:0] \address$17 ;
  input [3:0] endpoint;
  wire [3:0] endpoint;
  wire [3:0] \endpoint$18 ;
  output first;
  wire first;
  wire \first$11 ;
  wire \first$12 ;
  input [10:0] frame;
  wire [10:0] frame;
  wire [10:0] \frame$19 ;
  input is_in;
  wire is_in;
  input is_out;
  wire is_out;
  wire \is_out$21 ;
  input is_ping;
  wire is_ping;
  wire \is_ping$23 ;
  input is_setup;
  wire is_setup;
  wire \is_setup$22 ;
  output last;
  wire last;
  wire \last$13 ;
  input nak;
  wire nak;
  output \nak$2 ;
  wire \nak$2 ;
  wire \nak$28 ;
  input new_frame;
  wire new_frame;
  wire \new_frame$20 ;
  input new_token;
  wire new_token;
  input nyet;
  wire nyet;
  wire \nyet$26 ;
  wire \nyet$27 ;
  wire \nyet$30 ;
  output [7:0] payload;
  wire [7:0] payload;
  wire [7:0] \payload$14 ;
  input [3:0] pid;
  wire [3:0] pid;
  wire [3:0] \pid$16 ;
  input ready;
  wire ready;
  wire \ready$15 ;
  input ready_for_response;
  wire ready_for_response;
  input stall;
  wire stall;
  wire \stall$25 ;
  wire \stall$29 ;
  output \stall$3 ;
  wire \stall$3 ;
  wire tx_manager_ack;
  wire tx_manager_active;
  wire [1:0] tx_manager_data_pid;
  wire tx_manager_first;
  wire tx_manager_generate_zlps;
  wire tx_manager_is_in;
  wire tx_manager_last;
  wire \tx_manager_last$5 ;
  wire tx_manager_nak;
  wire tx_manager_new_token;
  wire [7:0] tx_manager_payload;
  wire [7:0] \tx_manager_payload$6 ;
  wire tx_manager_ready;
  wire \tx_manager_ready$7 ;
  wire tx_manager_ready_for_response;
  wire tx_manager_valid;
  wire \tx_manager_valid$4 ;
  output [1:0] tx_pid_toggle;
  wire [1:0] tx_pid_toggle;
  input usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  output valid;
  wire valid;
  wire \valid$10 ;
  assign \$8  = endpoint ==  2'h3;
  tx_manager tx_manager (
    .ack(tx_manager_ack),
    .active(tx_manager_active),
    .data_pid(tx_manager_data_pid),
    .first(tx_manager_first),
    .generate_zlps(1'h1),
    .is_in(tx_manager_is_in),
    .last(1'h0),
    .\last$2 (\tx_manager_last$5 ),
    .nak(tx_manager_nak),
    .new_token(tx_manager_new_token),
    .payload(8'h00),
    .\payload$3 (\tx_manager_payload$6 ),
    .ready(tx_manager_ready),
    .\ready$4 (\tx_manager_ready$7 ),
    .ready_for_response(tx_manager_ready_for_response),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst),
    .valid(1'h0),
    .\valid$1 (\tx_manager_valid$4 )
  );
  assign \valid$10  = 1'h0;
  assign \first$12  = 1'h0;
  assign \last$13  = 1'h0;
  assign \payload$14  = 8'h00;
  assign \ack$24  = 1'h0;
  assign \stall$25  = 1'h0;
  assign \nyet$27  = 1'h0;
  assign \nyet$30  = nyet;
  assign \stall$29  = stall;
  assign \nak$28  = nak;
  assign tx_manager_ack = ack;
  assign \nyet$26  = 1'h0;
  assign \stall$3  = 1'h0;
  assign \nak$2  = tx_manager_nak;
  assign \ack$1  = 1'h0;
  assign \is_ping$23  = is_ping;
  assign \is_setup$22  = is_setup;
  assign \is_out$21  = is_out;
  assign tx_manager_is_in = is_in;
  assign \new_frame$20  = new_frame;
  assign \frame$19  = frame;
  assign tx_manager_ready_for_response = ready_for_response;
  assign tx_manager_new_token = new_token;
  assign \endpoint$18  = endpoint;
  assign \address$17  = address;
  assign \pid$16  = pid;
  assign tx_pid_toggle = tx_manager_data_pid;
  assign \tx_manager_ready$7  = ready;
  assign payload = \tx_manager_payload$6 ;
  assign last = \tx_manager_last$5 ;
  assign first = tx_manager_first;
  assign valid = \tx_manager_valid$4 ;
  assign \ready$15  = tx_manager_ready;
  assign tx_manager_payload = 8'h00;
  assign tx_manager_last = 1'h0;
  assign \first$11  = 1'h0;
  assign tx_manager_valid = 1'h0;
  assign tx_manager_active = \$8 ;
  assign tx_manager_generate_zlps = 1'h1;
endmodule
module USBStreamInEndpoint_2831507112816(first, last, payload, ready, usb_rst, usb_clk, ack, nak, stall, nyet, pid, address, endpoint, new_token, ready_for_response, frame, new_frame, is_in, is_out, is_setup, is_ping
, \ack$1 , \nak$2 , \stall$3 , \valid$4 , tx_pid_toggle, \payload$5 , \first$6 , \last$7 , \ready$8 , valid);
  wire \$13 ;
  input ack;
  wire ack;
  output \ack$1 ;
  wire \ack$1 ;
  wire \ack$24 ;
  input [6:0] address;
  wire [6:0] address;
  wire [6:0] \address$17 ;
  input [3:0] endpoint;
  wire [3:0] endpoint;
  wire [3:0] \endpoint$18 ;
  input first;
  wire first;
  wire \first$15 ;
  output \first$6 ;
  wire \first$6 ;
  input [10:0] frame;
  wire [10:0] frame;
  wire [10:0] \frame$19 ;
  input is_in;
  wire is_in;
  input is_out;
  wire is_out;
  wire \is_out$21 ;
  input is_ping;
  wire is_ping;
  wire \is_ping$23 ;
  input is_setup;
  wire is_setup;
  wire \is_setup$22 ;
  input last;
  wire last;
  output \last$7 ;
  wire \last$7 ;
  input nak;
  wire nak;
  output \nak$2 ;
  wire \nak$2 ;
  wire \nak$28 ;
  input new_frame;
  wire new_frame;
  wire \new_frame$20 ;
  input new_token;
  wire new_token;
  input nyet;
  wire nyet;
  wire \nyet$26 ;
  wire \nyet$27 ;
  wire \nyet$30 ;
  input [7:0] payload;
  wire [7:0] payload;
  output [7:0] \payload$5 ;
  wire [7:0] \payload$5 ;
  input [3:0] pid;
  wire [3:0] pid;
  wire [3:0] \pid$16 ;
  output ready;
  wire ready;
  input \ready$8 ;
  wire \ready$8 ;
  input ready_for_response;
  wire ready_for_response;
  input stall;
  wire stall;
  wire \stall$25 ;
  wire \stall$29 ;
  output \stall$3 ;
  wire \stall$3 ;
  wire tx_manager_ack;
  wire tx_manager_active;
  wire [1:0] tx_manager_data_pid;
  wire tx_manager_first;
  wire tx_manager_generate_zlps;
  wire tx_manager_is_in;
  wire tx_manager_last;
  wire \tx_manager_last$10 ;
  wire tx_manager_nak;
  wire tx_manager_new_token;
  wire [7:0] tx_manager_payload;
  wire [7:0] \tx_manager_payload$11 ;
  wire tx_manager_ready;
  wire \tx_manager_ready$12 ;
  wire tx_manager_ready_for_response;
  wire tx_manager_valid;
  wire \tx_manager_valid$9 ;
  output [1:0] tx_pid_toggle;
  wire [1:0] tx_pid_toggle;
  input usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  input valid;
  wire valid;
  output \valid$4 ;
  wire \valid$4 ;
  assign \$13  = endpoint ==  3'h4;
  \tx_manager$5  tx_manager (
    .ack(tx_manager_ack),
    .active(tx_manager_active),
    .data_pid(tx_manager_data_pid),
    .first(tx_manager_first),
    .generate_zlps(1'h1),
    .is_in(tx_manager_is_in),
    .last(tx_manager_last),
    .\last$2 (\tx_manager_last$10 ),
    .nak(tx_manager_nak),
    .new_token(tx_manager_new_token),
    .payload(tx_manager_payload),
    .\payload$3 (\tx_manager_payload$11 ),
    .ready(tx_manager_ready),
    .\ready$4 (\tx_manager_ready$12 ),
    .ready_for_response(tx_manager_ready_for_response),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst),
    .valid(tx_manager_valid),
    .\valid$1 (\tx_manager_valid$9 )
  );
  assign \ack$24  = 1'h0;
  assign \stall$25  = 1'h0;
  assign \nyet$27  = 1'h0;
  assign \nyet$30  = nyet;
  assign \stall$29  = stall;
  assign \nak$28  = nak;
  assign tx_manager_ack = ack;
  assign \nyet$26  = 1'h0;
  assign \stall$3  = 1'h0;
  assign \nak$2  = tx_manager_nak;
  assign \ack$1  = 1'h0;
  assign \is_ping$23  = is_ping;
  assign \is_setup$22  = is_setup;
  assign \is_out$21  = is_out;
  assign tx_manager_is_in = is_in;
  assign \new_frame$20  = new_frame;
  assign \frame$19  = frame;
  assign tx_manager_ready_for_response = ready_for_response;
  assign tx_manager_new_token = new_token;
  assign \endpoint$18  = endpoint;
  assign \address$17  = address;
  assign \pid$16  = pid;
  assign tx_pid_toggle = tx_manager_data_pid;
  assign \tx_manager_ready$12  = \ready$8 ;
  assign \payload$5  = \tx_manager_payload$11 ;
  assign \last$7  = \tx_manager_last$10 ;
  assign \first$6  = tx_manager_first;
  assign \valid$4  = \tx_manager_valid$9 ;
  assign ready = tx_manager_ready;
  assign tx_manager_payload = payload;
  assign tx_manager_last = last;
  assign \first$15  = first;
  assign tx_manager_valid = valid;
  assign tx_manager_active = \$13 ;
  assign tx_manager_generate_zlps = 1'h1;
endmodule
module USBStreamOutEndpoint(first, last, payload, ready, usb_rst, usb_clk, endpoint, ready_for_response, is_out, is_ping, \valid$1 , next, \payload$2 , rx_complete, rx_ready_for_response, rx_invalid, rx_pid_toggle, ack, nak, valid);
  reg \$auto$verilog_backend.cc:2083:dump_module$5  = 0;
  wire \$10 ;
  wire \$100 ;
  wire \$102 ;
  wire \$104 ;
  wire \$106 ;
  wire \$108 ;
  wire \$110 ;
  wire \$112 ;
  wire \$114 ;
  wire \$116 ;
  wire \$117 ;
  wire \$12 ;
  wire \$120 ;
  wire \$122 ;
  wire \$124 ;
  wire \$126 ;
  wire \$128 ;
  wire \$130 ;
  wire \$132 ;
  wire \$134 ;
  wire \$135 ;
  wire \$137 ;
  wire \$139 ;
  wire \$14 ;
  wire \$141 ;
  wire \$143 ;
  wire \$144 ;
  wire \$146 ;
  wire \$148 ;
  wire \$150 ;
  wire \$152 ;
  wire \$154 ;
  wire \$156 ;
  wire \$159 ;
  wire \$16 ;
  wire \$161 ;
  wire \$163 ;
  wire \$166 ;
  wire \$168 ;
  wire \$169 ;
  wire \$171 ;
  wire \$173 ;
  wire \$174 ;
  wire \$177 ;
  wire \$18 ;
  wire \$180 ;
  wire \$182 ;
  wire \$184 ;
  wire \$186 ;
  wire \$188 ;
  wire \$189 ;
  wire \$192 ;
  wire \$194 ;
  wire \$196 ;
  wire [9:0] \$198 ;
  wire [9:0] \$199 ;
  wire \$20 ;
  wire \$201 ;
  wire \$203 ;
  wire \$205 ;
  wire \$207 ;
  wire \$209 ;
  wire \$211 ;
  wire \$213 ;
  wire \$215 ;
  wire \$217 ;
  wire \$219 ;
  wire \$22 ;
  wire \$221 ;
  wire \$223 ;
  wire \$225 ;
  wire \$227 ;
  wire \$229 ;
  wire \$231 ;
  wire \$233 ;
  wire \$235 ;
  wire \$237 ;
  wire \$239 ;
  wire \$24 ;
  wire \$241 ;
  wire \$243 ;
  wire \$245 ;
  wire \$247 ;
  wire \$249 ;
  wire \$251 ;
  wire \$252 ;
  wire \$254 ;
  wire \$256 ;
  wire \$258 ;
  wire \$26 ;
  wire \$260 ;
  wire \$262 ;
  wire \$264 ;
  wire \$267 ;
  wire \$269 ;
  wire \$271 ;
  wire \$273 ;
  wire \$275 ;
  wire \$28 ;
  wire \$30 ;
  wire \$32 ;
  wire \$34 ;
  wire \$36 ;
  wire \$38 ;
  wire \$40 ;
  wire \$42 ;
  wire \$44 ;
  wire \$46 ;
  wire \$48 ;
  wire \$50 ;
  wire \$52 ;
  wire \$54 ;
  wire \$56 ;
  wire \$58 ;
  wire \$6 ;
  wire \$60 ;
  wire \$62 ;
  wire \$64 ;
  wire \$66 ;
  wire \$68 ;
  wire \$69 ;
  wire \$7 ;
  wire \$71 ;
  wire \$73 ;
  wire \$75 ;
  wire \$77 ;
  wire \$79 ;
  wire \$81 ;
  wire \$84 ;
  wire \$86 ;
  wire \$88 ;
  wire \$90 ;
  wire \$92 ;
  wire \$94 ;
  wire \$96 ;
  wire \$98 ;
  output ack;
  wire ack;
  wire boundary_detector_complete_in;
  wire boundary_detector_complete_out;
  wire boundary_detector_first;
  wire boundary_detector_invalid_in;
  wire boundary_detector_invalid_out;
  wire boundary_detector_last;
  wire boundary_detector_next;
  wire \boundary_detector_next$4 ;
  wire [7:0] boundary_detector_payload;
  wire [7:0] \boundary_detector_payload$3 ;
  wire boundary_detector_valid;
  wire \boundary_detector_valid$5 ;
  input [3:0] endpoint;
  wire [3:0] endpoint;
  reg expected_data_toggle = 1'h0;
  reg \expected_data_toggle$next ;
  wire fifo_empty;
  wire fifo_full;
  wire fifo_read_commit;
  wire [9:0] fifo_read_data;
  wire fifo_read_en;
  wire [9:0] fifo_space_available;
  wire fifo_write_commit;
  wire [9:0] fifo_write_data;
  wire fifo_write_discard;
  wire fifo_write_en;
  output first;
  wire first;
  input is_out;
  wire is_out;
  input is_ping;
  wire is_ping;
  output last;
  wire last;
  output nak;
  wire nak;
  input next;
  wire next;
  reg overflow = 1'h0;
  reg \overflow$next ;
  output [7:0] payload;
  wire [7:0] payload;
  input [7:0] \payload$2 ;
  wire [7:0] \payload$2 ;
  input ready;
  wire ready;
  input ready_for_response;
  wire ready_for_response;
  reg [8:0] rx_cnt = 9'h000;
  reg [8:0] \rx_cnt$next ;
  input rx_complete;
  wire rx_complete;
  input rx_invalid;
  wire rx_invalid;
  input [1:0] rx_pid_toggle;
  wire [1:0] rx_pid_toggle;
  input rx_ready_for_response;
  wire rx_ready_for_response;
  reg transfer_active = 1'h0;
  reg \transfer_active$next ;
  input usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  output valid;
  wire valid;
  input \valid$1 ;
  wire \valid$1 ;
  assign \$100  = \$96  &  \$98 ;
  assign \$102  = \$90  |  \$100 ;
  assign \$104  = endpoint ==  3'h4;
  assign \$106  = \$104  &  is_out;
  assign \$108  = \$106  &  is_out;
  assign \$10  = boundary_detector_last &  \$6 ;
  assign \$110  = \$108  &  rx_ready_for_response;
  assign \$112  = endpoint ==  3'h4;
  assign \$114  = \$112  &  is_out;
  assign \$117  = rx_pid_toggle ==  expected_data_toggle;
  assign \$116  = ~  \$117 ;
  assign \$120  = \$114  &  \$116 ;
  assign \$122  = \$110  &  \$120 ;
  assign \$124  = \$102  |  \$122 ;
  assign \$126  = endpoint ==  3'h4;
  assign \$128  = \$126  &  is_out;
  assign \$12  = ~  transfer_active;
  assign \$130  = \$128  &  is_out;
  assign \$132  = \$130  &  rx_ready_for_response;
  assign \$135  = endpoint ==  3'h4;
  assign \$137  = \$135  &  is_out;
  assign \$139  = rx_pid_toggle ==  expected_data_toggle;
  assign \$141  = \$137  &  \$139 ;
  assign \$144  = endpoint ==  3'h4;
  assign \$146  = \$144  &  is_out;
  assign \$148  = rx_pid_toggle ==  expected_data_toggle;
  assign \$14  = boundary_detector_first &  \$12 ;
  assign \$150  = \$146  &  \$148 ;
  assign \$152  = \$150  &  \boundary_detector_next$4 ;
  assign \$154  = \$152  &  \boundary_detector_valid$5 ;
  assign \$156  = \$154  &  fifo_full;
  assign \$143  = ~  \$156 ;
  assign \$159  = \$141  &  \$143 ;
  assign \$161  = ~  overflow;
  assign \$163  = \$159  &  \$161 ;
  assign \$134  = ~  \$163 ;
  assign \$166  = \$132  &  \$134 ;
  assign \$16  = endpoint ==  3'h4;
  assign \$169  = endpoint ==  3'h4;
  assign \$171  = \$169  &  is_out;
  assign \$174  = rx_pid_toggle ==  expected_data_toggle;
  assign \$173  = ~  \$174 ;
  assign \$177  = \$171  &  \$173 ;
  assign \$168  = ~  \$177 ;
  assign \$180  = \$166  &  \$168 ;
  assign \$182  = endpoint ==  3'h4;
  assign \$184  = \$182  &  is_ping;
  assign \$186  = \$184  &  ready_for_response;
  assign \$18  = \$16  &  is_out;
  assign \$189  = fifo_space_available >=  10'h200;
  assign \$188  = ~  \$189 ;
  assign \$192  = \$186  &  \$188 ;
  assign \$194  = \$180  |  \$192 ;
  assign \$196  = ~  fifo_empty;
  assign \$199  = rx_cnt +  1'h1;
  assign \$201  = endpoint ==  3'h4;
  assign \$203  = \$201  &  is_out;
  assign \$205  = rx_pid_toggle ==  expected_data_toggle;
  assign \$207  = \$203  &  \$205 ;
  assign \$20  = rx_pid_toggle ==  expected_data_toggle;
  assign \$209  = \$207  &  \boundary_detector_next$4 ;
  assign \$211  = \$209  &  \boundary_detector_valid$5 ;
  assign \$213  = \$211  &  fifo_full;
  assign \$215  = fifo_write_commit |  fifo_write_discard;
  assign \$217  = rx_cnt ==  9'h1ff;
  assign \$219  = endpoint ==  3'h4;
  assign \$221  = \$219  &  is_out;
  assign \$223  = rx_pid_toggle ==  expected_data_toggle;
  assign \$225  = \$221  &  \$223 ;
  assign \$227  = \$225  &  \boundary_detector_next$4 ;
  assign \$22  = \$18  &  \$20 ;
  assign \$229  = \$227  &  \boundary_detector_valid$5 ;
  assign \$231  = \$229  &  fifo_full;
  assign \$233  = fifo_write_commit |  fifo_write_discard;
  assign \$235  = endpoint ==  3'h4;
  assign \$237  = \$235  &  is_out;
  assign \$239  = \$237  &  is_out;
  assign \$241  = \$239  &  rx_ready_for_response;
  assign \$243  = endpoint ==  3'h4;
  assign \$245  = \$243  &  is_out;
  assign \$247  = rx_pid_toggle ==  expected_data_toggle;
  assign \$24  = \$22  &  \boundary_detector_next$4 ;
  assign \$249  = \$245  &  \$247 ;
  assign \$252  = endpoint ==  3'h4;
  assign \$254  = \$252  &  is_out;
  assign \$256  = rx_pid_toggle ==  expected_data_toggle;
  assign \$258  = \$254  &  \$256 ;
  assign \$260  = \$258  &  \boundary_detector_next$4 ;
  assign \$262  = \$260  &  \boundary_detector_valid$5 ;
  assign \$264  = \$262  &  fifo_full;
  assign \$251  = ~  \$264 ;
  assign \$267  = \$249  &  \$251 ;
  assign \$26  = \$24  &  \boundary_detector_valid$5 ;
  assign \$269  = ~  overflow;
  assign \$271  = \$267  &  \$269 ;
  assign \$273  = \$241  &  \$271 ;
  assign \$275  = ~  expected_data_toggle;
  always @(posedge usb_clk)
    rx_cnt <= \rx_cnt$next ;
  always @(posedge usb_clk)
    transfer_active <= \transfer_active$next ;
  always @(posedge usb_clk)
    overflow <= \overflow$next ;
  always @(posedge usb_clk)
    expected_data_toggle <= \expected_data_toggle$next ;
  assign \$28  = ~  fifo_full;
  assign \$30  = \$26  &  \$28 ;
  assign \$32  = endpoint ==  3'h4;
  assign \$34  = \$32  &  is_out;
  assign \$36  = \$34  &  boundary_detector_complete_out;
  assign \$38  = ~  overflow;
  assign \$40  = \$36  &  \$38 ;
  assign \$42  = endpoint ==  3'h4;
  assign \$44  = \$42  &  is_out;
  assign \$46  = boundary_detector_complete_out &  overflow;
  assign \$48  = boundary_detector_invalid_out |  \$46 ;
  assign \$50  = \$44  &  \$48 ;
  assign \$52  = endpoint ==  3'h4;
  assign \$54  = \$52  &  is_out;
  assign \$56  = \$54  &  is_out;
  assign \$58  = \$56  &  rx_ready_for_response;
  assign \$60  = endpoint ==  3'h4;
  assign \$62  = \$60  &  is_out;
  assign \$64  = rx_pid_toggle ==  expected_data_toggle;
  assign \$66  = \$62  &  \$64 ;
  assign \$69  = endpoint ==  3'h4;
  assign \$71  = \$69  &  is_out;
  assign \$73  = rx_pid_toggle ==  expected_data_toggle;
  assign \$75  = \$71  &  \$73 ;
  assign \$77  = \$75  &  \boundary_detector_next$4 ;
  assign \$7  = rx_cnt ==  9'h1ff;
  assign \$79  = \$77  &  \boundary_detector_valid$5 ;
  assign \$81  = \$79  &  fifo_full;
  assign \$68  = ~  \$81 ;
  assign \$84  = \$66  &  \$68 ;
  assign \$86  = ~  overflow;
  assign \$88  = \$84  &  \$86 ;
  assign \$6  = ~  \$7 ;
  assign \$90  = \$58  &  \$88 ;
  assign \$92  = endpoint ==  3'h4;
  assign \$94  = \$92  &  is_ping;
  assign \$96  = \$94  &  ready_for_response;
  assign \$98  = fifo_space_available >=  10'h200;
  boundary_detector boundary_detector (
    .complete_in(boundary_detector_complete_in),
    .complete_out(boundary_detector_complete_out),
    .first(boundary_detector_first),
    .invalid_in(boundary_detector_invalid_in),
    .invalid_out(boundary_detector_invalid_out),
    .last(boundary_detector_last),
    .next(boundary_detector_next),
    .\next$2 (\boundary_detector_next$4 ),
    .payload(boundary_detector_payload),
    .\payload$1 (\boundary_detector_payload$3 ),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst),
    .valid(boundary_detector_valid),
    .\valid$3 (\boundary_detector_valid$5 )
  );
  fifo fifo (
    .empty(fifo_empty),
    .full(fifo_full),
    .read_commit(1'h1),
    .read_data(fifo_read_data),
    .read_en(fifo_read_en),
    .space_available(fifo_space_available),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst),
    .write_commit(fifo_write_commit),
    .write_data(fifo_write_data),
    .write_discard(fifo_write_discard),
    .write_en(fifo_write_en)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \rx_cnt$next  = rx_cnt;
    casez (fifo_write_en)
      1'h1:
          \rx_cnt$next  = \$199 [8:0];
    endcase
    casez ({ \$215 , \$213  })
      2'b?1:
          ;
      2'b1?:
          \rx_cnt$next  = 9'h000;
    endcase
    casez (usb_rst)
      1'h1:
          \rx_cnt$next  = 9'h000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \transfer_active$next  = transfer_active;
    casez (fifo_write_en)
      1'h1:
          casez (boundary_detector_last)
            1'h1:
                \transfer_active$next  = \$217 ;
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \transfer_active$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \overflow$next  = overflow;
    casez ({ \$233 , \$231  })
      2'b?1:
          \overflow$next  = 1'h1;
      2'b1?:
          \overflow$next  = 1'h0;
    endcase
    casez (usb_rst)
      1'h1:
          \overflow$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \expected_data_toggle$next  = expected_data_toggle;
    casez (\$273 )
      1'h1:
          \expected_data_toggle$next  = \$275 ;
    endcase
    casez (usb_rst)
      1'h1:
          \expected_data_toggle$next  = 1'h0;
    endcase
  end
  assign \$198  = \$199 ;
  assign fifo_read_commit = 1'h1;
  assign fifo_read_en = ready;
  assign first = fifo_read_data[9];
  assign last = fifo_read_data[8];
  assign payload = fifo_read_data[7:0];
  assign valid = \$196 ;
  assign nak = \$194 ;
  assign ack = \$124 ;
  assign fifo_write_discard = \$50 ;
  assign fifo_write_commit = \$40 ;
  assign fifo_write_en = \$30 ;
  assign fifo_write_data[9] = \$14 ;
  assign fifo_write_data[8] = \$10 ;
  assign fifo_write_data[7:0] = \boundary_detector_payload$3 ;
  assign boundary_detector_invalid_in = rx_invalid;
  assign boundary_detector_complete_in = rx_complete;
  assign boundary_detector_payload = \payload$2 ;
  assign boundary_detector_next = next;
  assign boundary_detector_valid = \valid$1 ;
endmodule
module boundary_detector(usb_clk, valid, next, payload, complete_in, invalid_in, \payload$1 , last, first, \next$2 , \valid$3 , complete_out, invalid_out, usb_rst);
  reg \$auto$verilog_backend.cc:2083:dump_module$6  = 0;
  wire \$10 ;
  wire \$12 ;
  wire \$14 ;
  wire \$16 ;
  wire \$18 ;
  wire \$20 ;
  wire \$22 ;
  wire \$24 ;
  wire \$26 ;
  wire \$28 ;
  wire \$30 ;
  wire \$32 ;
  wire \$4 ;
  wire \$6 ;
  wire \$8 ;
  reg [7:0] buffered_byte = 8'h00;
  reg [7:0] \buffered_byte$next ;
  reg buffered_complete = 1'h0;
  reg \buffered_complete$next ;
  reg buffered_invalid = 1'h0;
  reg \buffered_invalid$next ;
  input complete_in;
  wire complete_in;
  output complete_out;
  reg complete_out = 1'h0;
  reg \complete_out$next ;
  output first;
  reg first = 1'h0;
  reg \first$next ;
  reg [1:0] fsm_state = 2'h0;
  reg [1:0] \fsm_state$next ;
  input invalid_in;
  wire invalid_in;
  output invalid_out;
  reg invalid_out = 1'h0;
  reg \invalid_out$next ;
  reg is_first_byte = 1'h0;
  reg \is_first_byte$next ;
  output last;
  reg last = 1'h0;
  reg \last$next ;
  input next;
  wire next;
  output \next$2 ;
  reg \next$2  = 1'h0;
  reg \next$2$next ;
  input [7:0] payload;
  wire [7:0] payload;
  output [7:0] \payload$1 ;
  reg [7:0] \payload$1  = 8'h00;
  reg [7:0] \payload$1$next ;
  input usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  input valid;
  wire valid;
  output \valid$3 ;
  reg \valid$3  = 1'h0;
  reg \valid$3$next ;
  assign \$10  = valid &  next;
  assign \$12  = ~  valid;
  assign \$14  = buffered_complete |  complete_in;
  assign \$16  = buffered_invalid |  invalid_in;
  assign \$18  = valid &  next;
  assign \$20  = valid &  next;
  assign \$22  = valid &  next;
  assign \$24  = valid &  next;
  assign \$26  = valid &  next;
  assign \$28  = ~  valid;
  assign \$30  = valid &  next;
  assign \$32  = ~  valid;
  always @(posedge usb_clk)
    \valid$3  <= \valid$3$next ;
  always @(posedge usb_clk)
    first <= \first$next ;
  always @(posedge usb_clk)
    last <= \last$next ;
  always @(posedge usb_clk)
    \next$2  <= \next$2$next ;
  always @(posedge usb_clk)
    buffered_complete <= \buffered_complete$next ;
  always @(posedge usb_clk)
    buffered_invalid <= \buffered_invalid$next ;
  always @(posedge usb_clk)
    complete_out <= \complete_out$next ;
  always @(posedge usb_clk)
    invalid_out <= \invalid_out$next ;
  always @(posedge usb_clk)
    buffered_byte <= \buffered_byte$next ;
  always @(posedge usb_clk)
    is_first_byte <= \is_first_byte$next ;
  always @(posedge usb_clk)
    fsm_state <= \fsm_state$next ;
  always @(posedge usb_clk)
    \payload$1  <= \payload$1$next ;
  assign \$4  = valid &  next;
  assign \$6  = ~  valid;
  assign \$8  = ~  valid;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$6 ) begin end
    \valid$3$next  = \valid$3 ;
    casez (fsm_state)
      2'h0:
          \valid$3$next  = 1'h0;
      2'h1:
          \valid$3$next  = 1'h1;
    endcase
    casez (usb_rst)
      1'h1:
          \valid$3$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$6 ) begin end
    \first$next  = first;
    casez (fsm_state)
      2'h0:
          \first$next  = 1'h0;
      2'h1:
        begin
          casez (\$4 )
            1'h1:
                \first$next  = is_first_byte;
          endcase
          casez (\$6 )
            1'h1:
                \first$next  = is_first_byte;
          endcase
        end
      2'h2:
          \first$next  = 1'h0;
    endcase
    casez (usb_rst)
      1'h1:
          \first$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$6 ) begin end
    \fsm_state$next  = fsm_state;
    casez (fsm_state)
      2'h0:
          casez (\$26 )
            1'h1:
                \fsm_state$next  = 2'h1;
          endcase
      2'h1:
          casez (\$28 )
            1'h1:
                \fsm_state$next  = 2'h2;
          endcase
      2'h2:
          \fsm_state$next  = 2'h0;
    endcase
    casez (usb_rst)
      1'h1:
          \fsm_state$next  = 2'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$6 ) begin end
    \payload$1$next  = \payload$1 ;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
        begin
          casez (\$30 )
            1'h1:
                \payload$1$next  = buffered_byte;
          endcase
          casez (\$32 )
            1'h1:
                \payload$1$next  = buffered_byte;
          endcase
        end
    endcase
    casez (usb_rst)
      1'h1:
          \payload$1$next  = 8'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$6 ) begin end
    \last$next  = last;
    casez (fsm_state)
      2'h0:
          \last$next  = 1'h0;
      2'h1:
          casez (\$8 )
            1'h1:
                \last$next  = 1'h1;
          endcase
      2'h2:
          \last$next  = 1'h0;
    endcase
    casez (usb_rst)
      1'h1:
          \last$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$6 ) begin end
    \next$2$next  = \next$2 ;
    casez (fsm_state)
      2'h0:
          \next$2$next  = 1'h0;
      2'h1:
        begin
          \next$2$next  = 1'h0;
          casez (\$10 )
            1'h1:
                \next$2$next  = 1'h1;
          endcase
          casez (\$12 )
            1'h1:
                \next$2$next  = 1'h1;
          endcase
        end
      2'h2:
          \next$2$next  = 1'h0;
    endcase
    casez (usb_rst)
      1'h1:
          \next$2$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$6 ) begin end
    \buffered_complete$next  = buffered_complete;
    casez (fsm_state)
      2'h0:
          \buffered_complete$next  = 1'h0;
      2'h1:
          \buffered_complete$next  = \$14 ;
    endcase
    casez (usb_rst)
      1'h1:
          \buffered_complete$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$6 ) begin end
    \buffered_invalid$next  = buffered_invalid;
    casez (fsm_state)
      2'h0:
          \buffered_invalid$next  = 1'h0;
      2'h1:
          \buffered_invalid$next  = \$16 ;
    endcase
    casez (usb_rst)
      1'h1:
          \buffered_invalid$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$6 ) begin end
    \complete_out$next  = complete_out;
    casez (fsm_state)
      2'h0:
          \complete_out$next  = 1'h0;
      2'h1:
          ;
      2'h2:
          \complete_out$next  = buffered_complete;
    endcase
    casez (usb_rst)
      1'h1:
          \complete_out$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$6 ) begin end
    \invalid_out$next  = invalid_out;
    casez (fsm_state)
      2'h0:
          \invalid_out$next  = 1'h0;
      2'h1:
          ;
      2'h2:
          \invalid_out$next  = buffered_invalid;
    endcase
    casez (usb_rst)
      1'h1:
          \invalid_out$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$6 ) begin end
    \buffered_byte$next  = buffered_byte;
    casez (fsm_state)
      2'h0:
          casez (\$18 )
            1'h1:
                \buffered_byte$next  = payload;
          endcase
      2'h1:
          casez (\$20 )
            1'h1:
                \buffered_byte$next  = payload;
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \buffered_byte$next  = 8'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$6 ) begin end
    \is_first_byte$next  = is_first_byte;
    casez (fsm_state)
      2'h0:
          casez (\$22 )
            1'h1:
                \is_first_byte$next  = 1'h1;
          endcase
      2'h1:
          casez (\$24 )
            1'h1:
                \is_first_byte$next  = 1'h0;
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \is_first_byte$next  = 1'h0;
    endcase
  end
endmodule
module control_translator(usb_clk, busy, \busy$1 , bus_idle, xcvr_select, term_select, op_mode, suspend, id_pullup, dm_pulldown, dp_pulldown, chrg_vbus, dischrg_vbus, use_external_vbus_indicator, done, address, write_data, read_request, write_request, usb_rst);
  reg \$auto$verilog_backend.cc:2083:dump_module$7  = 0;
  wire \$10 ;
  wire \$12 ;
  wire \$14 ;
  wire \$16 ;
  wire \$18 ;
  wire \$2 ;
  wire \$20 ;
  wire \$22 ;
  wire \$24 ;
  wire \$26 ;
  wire \$28 ;
  wire \$30 ;
  wire \$32 ;
  wire \$34 ;
  wire \$36 ;
  wire \$38 ;
  wire \$4 ;
  wire \$40 ;
  wire \$42 ;
  wire \$6 ;
  wire \$8 ;
  output [5:0] address;
  reg [5:0] address;
  input bus_idle;
  wire bus_idle;
  input busy;
  wire busy;
  output \busy$1 ;
  reg \busy$1  = 1'h0;
  reg \busy$1$next ;
  input chrg_vbus;
  wire chrg_vbus;
  reg [7:0] current_register_value_04 = 8'h41;
  reg [7:0] \current_register_value_04$next ;
  reg [7:0] current_register_value_0a = 8'h06;
  reg [7:0] \current_register_value_0a$next ;
  input dischrg_vbus;
  wire dischrg_vbus;
  input dm_pulldown;
  wire dm_pulldown;
  input done;
  wire done;
  input dp_pulldown;
  wire dp_pulldown;
  input id_pullup;
  wire id_pullup;
  input [1:0] op_mode;
  wire [1:0] op_mode;
  output read_request;
  wire read_request;
  input suspend;
  wire suspend;
  input term_select;
  wire term_select;
  input usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  input use_external_vbus_indicator;
  wire use_external_vbus_indicator;
  output [7:0] write_data;
  reg [7:0] write_data;
  reg write_done_04;
  reg write_done_0a;
  output write_request;
  reg write_request;
  wire write_requested_04;
  wire write_requested_0a;
  reg [7:0] write_value_04 = 8'h00;
  reg [7:0] \write_value_04$next ;
  reg [7:0] write_value_0a = 8'h00;
  reg [7:0] \write_value_0a$next ;
  input [1:0] xcvr_select;
  wire [1:0] xcvr_select;
  assign \$10  = ~  suspend;
  assign \$12  = current_register_value_0a !=  { use_external_vbus_indicator, 2'h0, chrg_vbus, dischrg_vbus, dm_pulldown, dp_pulldown, id_pullup };
  assign \$14  = current_register_value_0a !=  { use_external_vbus_indicator, 2'h0, chrg_vbus, dischrg_vbus, dm_pulldown, dp_pulldown, id_pullup };
  assign \$16  = ~  done;
  assign \$18  = write_requested_04 &  \$16 ;
  assign \$20  = \$18  &  bus_idle;
  assign \$22  = ~  done;
  assign \$24  = write_requested_0a &  \$22 ;
  assign \$26  = \$24  &  bus_idle;
  assign \$28  = ~  done;
  assign \$2  = ~  suspend;
  assign \$30  = write_requested_04 &  \$28 ;
  assign \$32  = \$30  &  bus_idle;
  assign \$34  = \$32  |  busy;
  assign \$36  = ~  done;
  assign \$38  = write_requested_0a &  \$36 ;
  assign \$40  = \$38  &  bus_idle;
  assign \$42  = \$40  |  busy;
  always @(posedge usb_clk)
    current_register_value_04 <= \current_register_value_04$next ;
  always @(posedge usb_clk)
    write_value_04 <= \write_value_04$next ;
  always @(posedge usb_clk)
    current_register_value_0a <= \current_register_value_0a$next ;
  always @(posedge usb_clk)
    write_value_0a <= \write_value_0a$next ;
  always @(posedge usb_clk)
    \busy$1  <= \busy$1$next ;
  assign \$4  = current_register_value_04 !=  { 1'h0, \$2 , 1'h0, op_mode, term_select, xcvr_select };
  assign \$6  = ~  suspend;
  assign \$8  = current_register_value_04 !=  { 1'h0, \$6 , 1'h0, op_mode, term_select, xcvr_select };
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$7 ) begin end
    \current_register_value_04$next  = current_register_value_04;
    casez (write_done_04)
      1'h1:
          \current_register_value_04$next  = write_value_04;
    endcase
    casez (usb_rst)
      1'h1:
          \current_register_value_04$next  = 8'h41;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$7 ) begin end
    casez ({ write_requested_0a, write_requested_04 })
      2'b?1:
          \busy$1$next  = \$34 ;
      2'b1?:
          \busy$1$next  = \$42 ;
      default:
          \busy$1$next  = busy;
    endcase
    casez (usb_rst)
      1'h1:
          \busy$1$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$7 ) begin end
    write_done_0a = 1'h0;
    casez ({ write_requested_0a, write_requested_04 })
      2'b?1:
          ;
      2'b1?:
          write_done_0a = done;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$7 ) begin end
    \write_value_04$next  = write_value_04;
    casez (\$8 )
      1'h1:
          \write_value_04$next  = { 1'h0, \$10 , 1'h0, op_mode, term_select, xcvr_select };
    endcase
    casez (usb_rst)
      1'h1:
          \write_value_04$next  = 8'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$7 ) begin end
    \current_register_value_0a$next  = current_register_value_0a;
    casez (write_done_0a)
      1'h1:
          \current_register_value_0a$next  = write_value_0a;
    endcase
    casez (usb_rst)
      1'h1:
          \current_register_value_0a$next  = 8'h06;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$7 ) begin end
    \write_value_0a$next  = write_value_0a;
    casez (\$14 )
      1'h1:
          \write_value_0a$next  = { use_external_vbus_indicator, 2'h0, chrg_vbus, dischrg_vbus, dm_pulldown, dp_pulldown, id_pullup };
    endcase
    casez (usb_rst)
      1'h1:
          \write_value_0a$next  = 8'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$7 ) begin end
    write_done_04 = 1'h0;
    casez ({ write_requested_0a, write_requested_04 })
      2'b?1:
          write_done_04 = done;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$7 ) begin end
    address = 6'h00;
    casez ({ write_requested_0a, write_requested_04 })
      2'b?1:
          address = 6'h04;
      2'b1?:
          address = 6'h0a;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$7 ) begin end
    write_data = 8'h00;
    casez ({ write_requested_0a, write_requested_04 })
      2'b?1:
          write_data = write_value_04;
      2'b1?:
          write_data = write_value_0a;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$7 ) begin end
    casez ({ write_requested_0a, write_requested_04 })
      2'b?1:
          write_request = \$20 ;
      2'b1?:
          write_request = \$26 ;
      default:
          write_request = 1'h0;
    endcase
  end
  assign read_request = 1'h0;
  assign write_requested_0a = \$12 ;
  assign write_requested_04 = \$4 ;
endmodule
module data_crc(rx_valid, tx_valid, tx_data, usb_rst, usb_clk, start, crc, \start$1 , \crc$2 , \start$3 , \crc$4 , rx_data);
  reg \$auto$verilog_backend.cc:2083:dump_module$8  = 0;
  wire \$10 ;
  wire \$100 ;
  wire \$102 ;
  wire \$104 ;
  wire \$106 ;
  wire \$108 ;
  wire \$110 ;
  wire \$112 ;
  wire \$114 ;
  wire \$116 ;
  wire \$118 ;
  wire \$12 ;
  wire \$120 ;
  wire \$122 ;
  wire \$124 ;
  wire \$126 ;
  wire \$128 ;
  wire \$130 ;
  wire \$132 ;
  wire \$134 ;
  wire \$136 ;
  wire \$138 ;
  wire \$14 ;
  wire \$140 ;
  wire \$142 ;
  wire \$144 ;
  wire \$146 ;
  wire \$148 ;
  wire \$150 ;
  wire \$152 ;
  wire \$154 ;
  wire \$156 ;
  wire \$158 ;
  wire \$16 ;
  wire \$160 ;
  wire \$162 ;
  wire \$164 ;
  wire \$166 ;
  wire \$168 ;
  wire \$170 ;
  wire \$172 ;
  wire \$174 ;
  wire \$176 ;
  wire \$178 ;
  wire \$18 ;
  wire \$180 ;
  wire \$182 ;
  wire \$184 ;
  wire \$186 ;
  wire \$188 ;
  wire \$190 ;
  wire \$192 ;
  wire \$194 ;
  wire \$196 ;
  wire \$198 ;
  wire \$20 ;
  wire \$200 ;
  wire \$202 ;
  wire \$204 ;
  wire \$206 ;
  wire \$208 ;
  wire \$210 ;
  wire \$212 ;
  wire \$214 ;
  wire \$216 ;
  wire \$218 ;
  wire \$22 ;
  wire \$220 ;
  wire \$222 ;
  wire \$224 ;
  wire \$226 ;
  wire \$228 ;
  wire \$230 ;
  wire \$232 ;
  wire \$234 ;
  wire \$236 ;
  wire \$238 ;
  wire \$24 ;
  wire \$240 ;
  wire \$242 ;
  wire \$244 ;
  wire \$246 ;
  wire \$248 ;
  wire \$250 ;
  wire \$252 ;
  wire \$254 ;
  wire \$256 ;
  wire \$258 ;
  wire \$26 ;
  wire \$260 ;
  wire \$262 ;
  wire \$264 ;
  wire \$266 ;
  wire \$268 ;
  wire \$270 ;
  wire \$272 ;
  wire \$274 ;
  wire \$276 ;
  wire \$278 ;
  wire \$28 ;
  wire \$280 ;
  wire [15:0] \$282 ;
  wire \$30 ;
  wire \$32 ;
  wire \$34 ;
  wire \$36 ;
  wire \$38 ;
  wire \$40 ;
  wire \$42 ;
  wire \$44 ;
  wire \$46 ;
  wire \$48 ;
  wire \$50 ;
  wire \$52 ;
  wire \$54 ;
  wire \$56 ;
  wire \$58 ;
  wire \$6 ;
  wire \$60 ;
  wire \$62 ;
  wire \$64 ;
  wire \$66 ;
  wire \$68 ;
  wire \$70 ;
  wire \$72 ;
  wire \$74 ;
  wire \$76 ;
  wire \$78 ;
  wire \$8 ;
  wire \$80 ;
  wire \$82 ;
  wire \$84 ;
  wire \$86 ;
  wire \$88 ;
  wire \$90 ;
  wire \$92 ;
  wire \$94 ;
  wire \$96 ;
  wire \$98 ;
  output [15:0] crc;
  wire [15:0] crc;
  output [15:0] \crc$2 ;
  wire [15:0] \crc$2 ;
  output [15:0] \crc$4 ;
  wire [15:0] \crc$4 ;
  reg [15:0] \crc$5  = 16'hffff;
  reg [15:0] \crc$5$next ;
  wire [15:0] output_crc;
  input [7:0] rx_data;
  wire [7:0] rx_data;
  input rx_valid;
  wire rx_valid;
  input start;
  wire start;
  input \start$1 ;
  wire \start$1 ;
  input \start$3 ;
  wire \start$3 ;
  input [7:0] tx_data;
  wire [7:0] tx_data;
  input tx_valid;
  wire tx_valid;
  input usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  assign \$100  = \$96  ^  \$98 ;
  assign \$102  = rx_data[0] ^  rx_data[1];
  assign \$104  = \crc$5 [14] ^  \crc$5 [15];
  assign \$106  = \$102  ^  \$104 ;
  assign \$108  = \$106  ^  \crc$5 [0];
  assign \$10  = rx_data[0] ^  rx_data[1];
  assign \$110  = rx_data[0] ^  \crc$5 [1];
  assign \$112  = \$110  ^  \crc$5 [15];
  assign \$114  = rx_data[0] ^  rx_data[1];
  assign \$116  = \$114  ^  rx_data[2];
  assign \$118  = \$116  ^  rx_data[3];
  assign \$120  = \$118  ^  rx_data[4];
  assign \$122  = \$120  ^  rx_data[5];
  assign \$124  = \$122  ^  rx_data[6];
  assign \$126  = \$124  ^  rx_data[7];
  assign \$128  = \crc$5 [7] ^  \crc$5 [8];
  assign \$12  = \$10  ^  rx_data[2];
  assign \$130  = \$128  ^  \crc$5 [9];
  assign \$132  = \$130  ^  \crc$5 [10];
  assign \$134  = \$132  ^  \crc$5 [11];
  assign \$136  = \$134  ^  \crc$5 [12];
  assign \$138  = \$136  ^  \crc$5 [13];
  assign \$140  = \$138  ^  \crc$5 [14];
  assign \$142  = \$140  ^  \crc$5 [15];
  assign \$144  = \$126  ^  \$142 ;
  assign \$146  = tx_data[0] ^  tx_data[1];
  assign \$148  = \$146  ^  tx_data[2];
  assign \$14  = \$12  ^  rx_data[3];
  assign \$150  = \$148  ^  tx_data[3];
  assign \$152  = \$150  ^  tx_data[4];
  assign \$154  = \$152  ^  tx_data[5];
  assign \$156  = \$154  ^  tx_data[6];
  assign \$158  = \$156  ^  tx_data[7];
  assign \$160  = \crc$5 [8] ^  \crc$5 [9];
  assign \$162  = \$160  ^  \crc$5 [10];
  assign \$164  = \$162  ^  \crc$5 [11];
  assign \$166  = \$164  ^  \crc$5 [12];
  assign \$168  = \$166  ^  \crc$5 [13];
  assign \$16  = \$14  ^  rx_data[4];
  assign \$170  = \$168  ^  \crc$5 [14];
  assign \$172  = \$170  ^  \crc$5 [15];
  assign \$174  = \$158  ^  \$172 ;
  assign \$176  = tx_data[0] ^  tx_data[1];
  assign \$178  = \$176  ^  tx_data[2];
  assign \$180  = \$178  ^  tx_data[3];
  assign \$182  = \$180  ^  tx_data[4];
  assign \$184  = \$182  ^  tx_data[5];
  assign \$186  = \$184  ^  tx_data[6];
  assign \$188  = \crc$5 [9] ^  \crc$5 [10];
  assign \$18  = \$16  ^  rx_data[5];
  assign \$190  = \$188  ^  \crc$5 [11];
  assign \$192  = \$190  ^  \crc$5 [12];
  assign \$194  = \$192  ^  \crc$5 [13];
  assign \$196  = \$194  ^  \crc$5 [14];
  assign \$198  = \$196  ^  \crc$5 [15];
  assign \$200  = \$186  ^  \$198 ;
  assign \$202  = tx_data[6] ^  tx_data[7];
  assign \$204  = \crc$5 [8] ^  \crc$5 [9];
  assign \$206  = \$202  ^  \$204 ;
  assign \$208  = tx_data[5] ^  tx_data[6];
  assign \$20  = \$18  ^  rx_data[6];
  assign \$210  = \crc$5 [9] ^  \crc$5 [10];
  assign \$212  = \$208  ^  \$210 ;
  assign \$214  = tx_data[4] ^  tx_data[5];
  assign \$216  = \crc$5 [10] ^  \crc$5 [11];
  assign \$218  = \$214  ^  \$216 ;
  assign \$220  = tx_data[3] ^  tx_data[4];
  assign \$222  = \crc$5 [11] ^  \crc$5 [12];
  assign \$224  = \$220  ^  \$222 ;
  assign \$226  = tx_data[2] ^  tx_data[3];
  assign \$228  = \crc$5 [12] ^  \crc$5 [13];
  assign \$22  = \$20  ^  rx_data[7];
  assign \$230  = \$226  ^  \$228 ;
  assign \$232  = tx_data[1] ^  tx_data[2];
  assign \$234  = \crc$5 [13] ^  \crc$5 [14];
  assign \$236  = \$232  ^  \$234 ;
  assign \$238  = tx_data[0] ^  tx_data[1];
  assign \$240  = \crc$5 [14] ^  \crc$5 [15];
  assign \$242  = \$238  ^  \$240 ;
  assign \$244  = \$242  ^  \crc$5 [0];
  assign \$246  = tx_data[0] ^  \crc$5 [1];
  assign \$248  = \$246  ^  \crc$5 [15];
  assign \$24  = \crc$5 [8] ^  \crc$5 [9];
  assign \$250  = tx_data[0] ^  tx_data[1];
  assign \$252  = \$250  ^  tx_data[2];
  assign \$254  = \$252  ^  tx_data[3];
  assign \$256  = \$254  ^  tx_data[4];
  assign \$258  = \$256  ^  tx_data[5];
  assign \$260  = \$258  ^  tx_data[6];
  assign \$262  = \$260  ^  tx_data[7];
  assign \$264  = \crc$5 [7] ^  \crc$5 [8];
  assign \$266  = \$264  ^  \crc$5 [9];
  assign \$268  = \$266  ^  \crc$5 [10];
  assign \$26  = \$24  ^  \crc$5 [10];
  assign \$270  = \$268  ^  \crc$5 [11];
  assign \$272  = \$270  ^  \crc$5 [12];
  assign \$274  = \$272  ^  \crc$5 [13];
  assign \$276  = \$274  ^  \crc$5 [14];
  assign \$278  = \$276  ^  \crc$5 [15];
  assign \$280  = \$262  ^  \$278 ;
  assign \$282  = ~  { \crc$5 [0], \crc$5 [1], \crc$5 [2], \crc$5 [3], \crc$5 [4], \crc$5 [5], \crc$5 [6], \crc$5 [7], \crc$5 [8], \crc$5 [9], \crc$5 [10], \crc$5 [11], \crc$5 [12], \crc$5 [13], \crc$5 [14], \crc$5 [15] };
  always @(posedge usb_clk)
    \crc$5  <= \crc$5$next ;
  assign \$28  = \$26  ^  \crc$5 [11];
  assign \$30  = \$28  ^  \crc$5 [12];
  assign \$32  = \$30  ^  \crc$5 [13];
  assign \$34  = \$32  ^  \crc$5 [14];
  assign \$36  = \$34  ^  \crc$5 [15];
  assign \$38  = \$22  ^  \$36 ;
  assign \$40  = rx_data[0] ^  rx_data[1];
  assign \$42  = \$40  ^  rx_data[2];
  assign \$44  = \$42  ^  rx_data[3];
  assign \$46  = \$44  ^  rx_data[4];
  assign \$48  = \$46  ^  rx_data[5];
  assign \$50  = \$48  ^  rx_data[6];
  assign \$52  = \crc$5 [9] ^  \crc$5 [10];
  assign \$54  = \$52  ^  \crc$5 [11];
  assign \$56  = \$54  ^  \crc$5 [12];
  assign \$58  = \$56  ^  \crc$5 [13];
  assign \$60  = \$58  ^  \crc$5 [14];
  assign \$62  = \$60  ^  \crc$5 [15];
  assign \$64  = \$50  ^  \$62 ;
  assign \$66  = rx_data[6] ^  rx_data[7];
  assign \$68  = \crc$5 [8] ^  \crc$5 [9];
  assign \$6  = start |  \start$1 ;
  assign \$70  = \$66  ^  \$68 ;
  assign \$72  = rx_data[5] ^  rx_data[6];
  assign \$74  = \crc$5 [9] ^  \crc$5 [10];
  assign \$76  = \$72  ^  \$74 ;
  assign \$78  = rx_data[4] ^  rx_data[5];
  assign \$80  = \crc$5 [10] ^  \crc$5 [11];
  assign \$82  = \$78  ^  \$80 ;
  assign \$84  = rx_data[3] ^  rx_data[4];
  assign \$86  = \crc$5 [11] ^  \crc$5 [12];
  assign \$88  = \$84  ^  \$86 ;
  assign \$8  = \$6  |  \start$3 ;
  assign \$90  = rx_data[2] ^  rx_data[3];
  assign \$92  = \crc$5 [12] ^  \crc$5 [13];
  assign \$94  = \$90  ^  \$92 ;
  assign \$96  = rx_data[1] ^  rx_data[2];
  assign \$98  = \crc$5 [13] ^  \crc$5 [14];
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$8 ) begin end
    \crc$5$next  = \crc$5 ;
    casez ({ tx_valid, rx_valid, \$8  })
      3'b??1:
          \crc$5$next  = 16'hffff;
      3'b?1?:
          \crc$5$next  = { \$144 , \crc$5 [6:2], \$112 , \$108 , \$100 , \$94 , \$88 , \$82 , \$76 , \$70 , \$64 , \$38  };
      3'b1??:
          \crc$5$next  = { \$280 , \crc$5 [6:2], \$248 , \$244 , \$236 , \$230 , \$224 , \$218 , \$212 , \$206 , \$200 , \$174  };
    endcase
    casez (usb_rst)
      1'h1:
          \crc$5$next  = 16'hffff;
    endcase
  end
  assign \crc$4  = output_crc;
  assign \crc$2  = output_crc;
  assign crc = output_crc;
  assign output_crc = \$282 ;
endmodule
module data_handler(rx_valid, usb_rst, usb_clk, rx_active, start, crc, new_packet, length, packet_0, packet_1, packet_2, packet_3, packet_4, packet_5, packet_6, packet_7, rx_data);
  reg \$auto$verilog_backend.cc:2083:dump_module$9  = 0;
  wire \$1 ;
  wire \$100 ;
  wire \$102 ;
  wire \$104 ;
  wire \$106 ;
  wire \$11 ;
  wire \$13 ;
  wire \$15 ;
  wire \$17 ;
  wire \$19 ;
  wire \$21 ;
  wire \$23 ;
  wire [3:0] \$25 ;
  wire \$27 ;
  wire \$29 ;
  wire \$3 ;
  wire \$31 ;
  wire \$33 ;
  wire [3:0] \$35 ;
  wire \$37 ;
  wire \$39 ;
  wire \$41 ;
  wire \$43 ;
  wire [4:0] \$45 ;
  wire [4:0] \$46 ;
  wire \$5 ;
  wire \$57 ;
  wire \$59 ;
  wire \$61 ;
  wire \$63 ;
  wire \$65 ;
  wire \$67 ;
  wire \$69 ;
  wire [3:0] \$7 ;
  wire \$71 ;
  wire [4:0] \$73 ;
  wire [4:0] \$74 ;
  wire \$76 ;
  wire \$78 ;
  wire \$80 ;
  wire \$82 ;
  wire \$84 ;
  wire \$86 ;
  wire \$88 ;
  wire \$9 ;
  wire \$90 ;
  wire \$92 ;
  wire \$94 ;
  wire \$96 ;
  wire \$98 ;
  reg [7:0] \$signal  = 8'h00;
  reg [7:0] \$signal$48  = 8'h00;
  reg [7:0] \$signal$48$next ;
  reg [7:0] \$signal$49  = 8'h00;
  reg [7:0] \$signal$49$next ;
  reg [7:0] \$signal$50  = 8'h00;
  reg [7:0] \$signal$50$next ;
  reg [7:0] \$signal$51  = 8'h00;
  reg [7:0] \$signal$51$next ;
  reg [7:0] \$signal$52  = 8'h00;
  reg [7:0] \$signal$52$next ;
  reg [7:0] \$signal$53  = 8'h00;
  reg [7:0] \$signal$53$next ;
  reg [7:0] \$signal$54  = 8'h00;
  reg [7:0] \$signal$54$next ;
  reg [7:0] \$signal$55  = 8'h00;
  reg [7:0] \$signal$55$next ;
  reg [7:0] \$signal$56  = 8'h00;
  reg [7:0] \$signal$56$next ;
  reg [7:0] \$signal$next ;
  reg [3:0] active_pid = 4'h0;
  reg [3:0] \active_pid$next ;
  input [15:0] crc;
  wire [15:0] crc;
  reg [1:0] fsm_state = 2'h0;
  reg [1:0] \fsm_state$next ;
  reg [15:0] last_byte_crc = 16'h0000;
  reg [15:0] \last_byte_crc$next ;
  reg [15:0] last_word = 16'h0000;
  reg [15:0] \last_word$next ;
  reg [15:0] last_word_crc = 16'h0000;
  reg [15:0] \last_word_crc$next ;
  output [3:0] length;
  reg [3:0] length = 4'h0;
  reg [3:0] \length$next ;
  output new_packet;
  reg new_packet = 1'h0;
  reg \new_packet$next ;
  output [7:0] packet_0;
  reg [7:0] packet_0 = 8'h00;
  reg [7:0] \packet_0$next ;
  output [7:0] packet_1;
  reg [7:0] packet_1 = 8'h00;
  reg [7:0] \packet_1$next ;
  output [7:0] packet_2;
  reg [7:0] packet_2 = 8'h00;
  reg [7:0] \packet_2$next ;
  output [7:0] packet_3;
  reg [7:0] packet_3 = 8'h00;
  reg [7:0] \packet_3$next ;
  output [7:0] packet_4;
  reg [7:0] packet_4 = 8'h00;
  reg [7:0] \packet_4$next ;
  output [7:0] packet_5;
  reg [7:0] packet_5 = 8'h00;
  reg [7:0] \packet_5$next ;
  output [7:0] packet_6;
  reg [7:0] packet_6 = 8'h00;
  reg [7:0] \packet_6$next ;
  output [7:0] packet_7;
  reg [7:0] packet_7 = 8'h00;
  reg [7:0] \packet_7$next ;
  reg [3:0] packet_id = 4'h0;
  reg [3:0] \packet_id$next ;
  reg [3:0] position_in_packet = 4'h0;
  reg [3:0] \position_in_packet$next ;
  input rx_active;
  wire rx_active;
  input [7:0] rx_data;
  wire [7:0] rx_data;
  input rx_valid;
  wire rx_valid;
  output start;
  reg start;
  input usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  assign \$9  = rx_data[3:0] ==  \$7 ;
  assign \$100  = ~  rx_active;
  assign \$102  = last_word_crc ==  last_word;
  assign \$104  = ~  rx_active;
  assign \$106  = last_word_crc ==  last_word;
  always @(posedge usb_clk)
    new_packet <= \new_packet$next ;
  always @(posedge usb_clk)
    fsm_state <= \fsm_state$next ;
  always @(posedge usb_clk)
    active_pid <= \active_pid$next ;
  always @(posedge usb_clk)
    position_in_packet <= \position_in_packet$next ;
  always @(posedge usb_clk)
    \$signal  <= \$signal$next ;
  always @(posedge usb_clk)
    \$signal$48  <= \$signal$48$next ;
  always @(posedge usb_clk)
    \$signal$49  <= \$signal$49$next ;
  always @(posedge usb_clk)
    \$signal$50  <= \$signal$50$next ;
  always @(posedge usb_clk)
    \$signal$51  <= \$signal$51$next ;
  always @(posedge usb_clk)
    \$signal$52  <= \$signal$52$next ;
  always @(posedge usb_clk)
    \$signal$53  <= \$signal$53$next ;
  always @(posedge usb_clk)
    \$signal$54  <= \$signal$54$next ;
  assign \$11  = rx_data[1:0] ==  2'h3;
  always @(posedge usb_clk)
    \$signal$55  <= \$signal$55$next ;
  always @(posedge usb_clk)
    \$signal$56  <= \$signal$56$next ;
  always @(posedge usb_clk)
    last_word <= \last_word$next ;
  always @(posedge usb_clk)
    last_word_crc <= \last_word_crc$next ;
  always @(posedge usb_clk)
    last_byte_crc <= \last_byte_crc$next ;
  always @(posedge usb_clk)
    packet_id <= \packet_id$next ;
  always @(posedge usb_clk)
    length <= \length$next ;
  always @(posedge usb_clk)
    packet_0 <= \packet_0$next ;
  always @(posedge usb_clk)
    packet_1 <= \packet_1$next ;
  always @(posedge usb_clk)
    packet_2 <= \packet_2$next ;
  always @(posedge usb_clk)
    packet_3 <= \packet_3$next ;
  always @(posedge usb_clk)
    packet_4 <= \packet_4$next ;
  always @(posedge usb_clk)
    packet_5 <= \packet_5$next ;
  always @(posedge usb_clk)
    packet_6 <= \packet_6$next ;
  always @(posedge usb_clk)
    packet_7 <= \packet_7$next ;
  assign \$13  = \$9  &  \$11 ;
  assign \$15  = position_in_packet >=  4'ha;
  assign \$17  = ~  rx_active;
  assign \$1  = ~  rx_active;
  assign \$19  = last_word_crc ==  last_word;
  assign \$21  = ~  rx_active;
  assign \$23  = ~  rx_active;
  assign \$25  = ~  rx_data[7:4];
  assign \$27  = rx_data[3:0] ==  \$25 ;
  assign \$29  = rx_data[1:0] ==  2'h3;
  assign \$31  = \$27  &  \$29 ;
  assign \$33  = ~  rx_active;
  assign \$35  = ~  rx_data[7:4];
  assign \$37  = rx_data[3:0] ==  \$35 ;
  assign \$3  = last_word_crc ==  last_word;
  assign \$39  = rx_data[1:0] ==  2'h3;
  assign \$41  = \$37  &  \$39 ;
  assign \$43  = position_in_packet >=  4'ha;
  assign \$46  = position_in_packet +  1'h1;
  assign \$57  = position_in_packet >=  4'ha;
  assign \$5  = ~  rx_active;
  assign \$59  = position_in_packet >=  4'ha;
  assign \$61  = position_in_packet >=  4'ha;
  assign \$63  = position_in_packet >=  4'ha;
  assign \$65  = ~  rx_active;
  assign \$67  = last_word_crc ==  last_word;
  assign \$69  = ~  rx_active;
  assign \$71  = last_word_crc ==  last_word;
  assign \$74  = position_in_packet -  2'h2;
  assign \$76  = ~  rx_active;
  assign \$78  = last_word_crc ==  last_word;
  assign \$7  = ~  rx_data[7:4];
  assign \$80  = ~  rx_active;
  assign \$82  = last_word_crc ==  last_word;
  assign \$84  = ~  rx_active;
  assign \$86  = last_word_crc ==  last_word;
  assign \$88  = ~  rx_active;
  assign \$90  = last_word_crc ==  last_word;
  assign \$92  = ~  rx_active;
  assign \$94  = last_word_crc ==  last_word;
  assign \$96  = ~  rx_active;
  assign \$98  = last_word_crc ==  last_word;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$9 ) begin end
    \new_packet$next  = 1'h0;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          ;
      2'h2:
          casez (\$1 )
            1'h1:
                casez (\$3 )
                  1'h1:
                      \new_packet$next  = 1'h1;
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \new_packet$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$9 ) begin end
    start = 1'h0;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          start = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$9 ) begin end
    \last_word$next  = last_word;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          ;
      2'h2:
          casez (rx_valid)
            1'h1:
                casez (\$59 )
                  1'h1:
                      ;
                  default:
                      \last_word$next  = { rx_data, last_word[15:8] };
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \last_word$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$9 ) begin end
    \last_word_crc$next  = last_word_crc;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          ;
      2'h2:
          casez (rx_valid)
            1'h1:
                casez (\$61 )
                  1'h1:
                      ;
                  default:
                      \last_word_crc$next  = last_byte_crc;
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \last_word_crc$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$9 ) begin end
    \last_byte_crc$next  = last_byte_crc;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          ;
      2'h2:
          casez (rx_valid)
            1'h1:
                casez (\$63 )
                  1'h1:
                      ;
                  default:
                      \last_byte_crc$next  = crc;
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \last_byte_crc$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$9 ) begin end
    \packet_id$next  = packet_id;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          ;
      2'h2:
          casez (\$65 )
            1'h1:
                casez (\$67 )
                  1'h1:
                      \packet_id$next  = active_pid;
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \packet_id$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$9 ) begin end
    \length$next  = length;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          ;
      2'h2:
          casez (\$69 )
            1'h1:
                casez (\$71 )
                  1'h1:
                      \length$next  = \$74 [3:0];
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \length$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$9 ) begin end
    \fsm_state$next  = fsm_state;
    casez (fsm_state)
      2'h0:
          casez (rx_active)
            1'h1:
                \fsm_state$next  = 2'h1;
          endcase
      2'h1:
          casez ({ rx_valid, \$5  })
            2'b?1:
                \fsm_state$next  = 2'h0;
            2'b1?:
                casez (\$13 )
                  1'h1:
                      \fsm_state$next  = 2'h2;
                  default:
                      \fsm_state$next  = 2'h3;
                endcase
          endcase
      2'h2:
        begin
          casez (rx_valid)
            1'h1:
                casez (\$15 )
                  1'h1:
                      \fsm_state$next  = 2'h3;
                endcase
          endcase
          casez (\$17 )
            1'h1:
                casez (\$19 )
                  1'h1:
                      \fsm_state$next  = 2'h0;
                endcase
          endcase
        end
      2'h3:
          casez (\$21 )
            1'h1:
                \fsm_state$next  = 2'h0;
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \fsm_state$next  = 2'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$9 ) begin end
    \packet_0$next  = packet_0;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          ;
      2'h2:
          casez (\$76 )
            1'h1:
                casez (\$78 )
                  1'h1:
                      \packet_0$next  = \$signal ;
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \packet_0$next  = 8'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$9 ) begin end
    \packet_1$next  = packet_1;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          ;
      2'h2:
          casez (\$80 )
            1'h1:
                casez (\$82 )
                  1'h1:
                      \packet_1$next  = \$signal$48 ;
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \packet_1$next  = 8'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$9 ) begin end
    \packet_2$next  = packet_2;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          ;
      2'h2:
          casez (\$84 )
            1'h1:
                casez (\$86 )
                  1'h1:
                      \packet_2$next  = \$signal$49 ;
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \packet_2$next  = 8'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$9 ) begin end
    \packet_3$next  = packet_3;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          ;
      2'h2:
          casez (\$88 )
            1'h1:
                casez (\$90 )
                  1'h1:
                      \packet_3$next  = \$signal$50 ;
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \packet_3$next  = 8'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$9 ) begin end
    \packet_4$next  = packet_4;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          ;
      2'h2:
          casez (\$92 )
            1'h1:
                casez (\$94 )
                  1'h1:
                      \packet_4$next  = \$signal$51 ;
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \packet_4$next  = 8'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$9 ) begin end
    \packet_5$next  = packet_5;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          ;
      2'h2:
          casez (\$96 )
            1'h1:
                casez (\$98 )
                  1'h1:
                      \packet_5$next  = \$signal$52 ;
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \packet_5$next  = 8'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$9 ) begin end
    \packet_6$next  = packet_6;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          ;
      2'h2:
          casez (\$100 )
            1'h1:
                casez (\$102 )
                  1'h1:
                      \packet_6$next  = \$signal$53 ;
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \packet_6$next  = 8'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$9 ) begin end
    \packet_7$next  = packet_7;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          ;
      2'h2:
          casez (\$104 )
            1'h1:
                casez (\$106 )
                  1'h1:
                      \packet_7$next  = \$signal$54 ;
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \packet_7$next  = 8'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$9 ) begin end
    \active_pid$next  = active_pid;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          casez ({ rx_valid, \$23  })
            2'b?1:
                ;
            2'b1?:
                casez (\$31 )
                  1'h1:
                      \active_pid$next  = rx_data[3:0];
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \active_pid$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$9 ) begin end
    \position_in_packet$next  = position_in_packet;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          casez ({ rx_valid, \$33  })
            2'b?1:
                ;
            2'b1?:
                casez (\$41 )
                  1'h1:
                      \position_in_packet$next  = 4'h0;
                endcase
          endcase
      2'h2:
          casez (rx_valid)
            1'h1:
                casez (\$43 )
                  1'h1:
                      ;
                  default:
                      \position_in_packet$next  = \$46 [3:0];
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \position_in_packet$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$9 ) begin end
    \$signal$next  = \$signal ;
    \$signal$48$next  = \$signal$48 ;
    \$signal$49$next  = \$signal$49 ;
    \$signal$50$next  = \$signal$50 ;
    \$signal$51$next  = \$signal$51 ;
    \$signal$52$next  = \$signal$52 ;
    \$signal$53$next  = \$signal$53 ;
    \$signal$54$next  = \$signal$54 ;
    \$signal$55$next  = \$signal$55 ;
    \$signal$56$next  = \$signal$56 ;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          ;
      2'h2:
          casez (rx_valid)
            1'h1:
                casez (\$57 )
                  1'h1:
                      ;
                  default:
                      casez (position_in_packet)
                        4'h0:
                            \$signal$next  = rx_data;
                        4'h1:
                            \$signal$48$next  = rx_data;
                        4'h2:
                            \$signal$49$next  = rx_data;
                        4'h3:
                            \$signal$50$next  = rx_data;
                        4'h4:
                            \$signal$51$next  = rx_data;
                        4'h5:
                            \$signal$52$next  = rx_data;
                        4'h6:
                            \$signal$53$next  = rx_data;
                        4'h7:
                            \$signal$54$next  = rx_data;
                        4'h8:
                            \$signal$55$next  = rx_data;
                        4'h?:
                            \$signal$56$next  = rx_data;
                      endcase
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
        begin
          \$signal$next  = 8'h00;
          \$signal$48$next  = 8'h00;
          \$signal$49$next  = 8'h00;
          \$signal$50$next  = 8'h00;
          \$signal$51$next  = 8'h00;
          \$signal$52$next  = 8'h00;
          \$signal$53$next  = 8'h00;
          \$signal$54$next  = 8'h00;
          \$signal$55$next  = 8'h00;
          \$signal$56$next  = 8'h00;
        end
    endcase
  end
  assign \$45  = \$46 ;
  assign \$73  = \$74 ;
endmodule
module encoder(o, i);
  reg \$auto$verilog_backend.cc:2083:dump_module$10  = 0;
  input [3:0] i;
  wire [3:0] i;
  reg n;
  output [1:0] o;
  reg [1:0] o;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$10 ) begin end
    o = 2'h0;
    casez (i)
      4'h1:
          o = 2'h0;
      4'h2:
          o = 2'h1;
      4'h4:
          o = 2'h2;
      4'h8:
          o = 2'h3;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$10 ) begin end
    n = 1'h0;
    casez (i)
      4'h1:
          ;
      4'h2:
          ;
      4'h4:
          ;
      4'h8:
          ;
      default:
          n = 1'h1;
    endcase
  end
endmodule
module \encoder$3 (o, i);
  reg \$auto$verilog_backend.cc:2083:dump_module$11  = 0;
  input [2:0] i;
  wire [2:0] i;
  reg n;
  output [1:0] o;
  reg [1:0] o;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$11 ) begin end
    o = 2'h0;
    casez (i)
      3'h1:
          o = 2'h0;
      3'h2:
          o = 2'h1;
      3'h4:
          o = 2'h2;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$11 ) begin end
    n = 1'h0;
    casez (i)
      3'h1:
          ;
      3'h2:
          ;
      3'h4:
          ;
      default:
          n = 1'h1;
    endcase
  end
endmodule
module \encoder$6 (o, i);
  reg \$auto$verilog_backend.cc:2083:dump_module$12  = 0;
  input [2:0] i;
  wire [2:0] i;
  reg n;
  output [1:0] o;
  reg [1:0] o;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$12 ) begin end
    o = 2'h0;
    casez (i)
      3'h1:
          o = 2'h0;
      3'h2:
          o = 2'h1;
      3'h4:
          o = 2'h2;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$12 ) begin end
    n = 1'h0;
    casez (i)
      3'h1:
          ;
      3'h2:
          ;
      3'h4:
          ;
      default:
          n = 1'h1;
    endcase
  end
endmodule
module endpoint_mux(address, endpoint, new_token, ready_for_response, frame, new_frame, is_in, is_out, is_setup, is_ping, ack, nak, stall, nyet, speed, active_config, active_address, valid, next, payload, rx_complete
, rx_invalid, rx_ready_for_response, rx_pid_toggle, \valid$1 , first, last, \payload$2 , ready, \ack$3 , \nak$4 , \stall$5 , tx_pid_toggle, address_changed, new_address, config_changed, new_config, usb_rst, usb_clk, start, crc, \start$6 
, tx_allowed, tx_timeout, rx_timeout, \crc$7 , \tx_allowed$8 , \tx_timeout$9 , \rx_timeout$10 , \ack$11 , \nak$12 , \stall$13 , \nyet$14 , \pid$15 , \address$16 , \endpoint$17 , \new_token$18 , \ready_for_response$19 , \frame$20 , \new_frame$21 , \is_in$22 , \is_out$23 , \is_setup$24 
, \is_ping$25 , \valid$26 , \next$27 , \payload$28 , \rx_ready_for_response$29 , \speed$30 , \active_config$31 , \ack$32 , \nak$33 , \stall$34 , \nyet$35 , \pid$36 , \address$37 , \endpoint$38 , \new_token$39 , \ready_for_response$40 , \frame$41 , \new_frame$42 , \is_in$43 , \is_out$44 , \is_setup$45 
, \is_ping$46 , \endpoint$47 , \ready_for_response$48 , \is_out$49 , \is_ping$50 , \valid$51 , \next$52 , \payload$53 , \rx_complete$54 , \rx_ready_for_response$55 , \rx_invalid$56 , \rx_pid_toggle$57 , \ack$58 , \nak$59 , \stall$60 , \nyet$61 , \pid$62 , \address$63 , \endpoint$64 , \new_token$65 , \ready_for_response$66 
, \frame$67 , \new_frame$68 , \is_in$69 , \is_out$70 , \is_setup$71 , \is_ping$72 , \address_changed$73 , \new_address$74 , \config_changed$75 , \new_config$76 , \ack$77 , \ack$78 , \ack$79 , \ack$80 , \nak$81 , \nak$82 , \nak$83 , \nak$84 , \stall$85 , \stall$86 , \stall$87 
, \start$88 , \start$89 , \valid$90 , \valid$91 , \valid$92 , \tx_pid_toggle$93 , \tx_pid_toggle$94 , \tx_pid_toggle$95 , \payload$96 , \payload$97 , \payload$98 , \first$99 , \first$100 , \first$101 , \last$102 , \last$103 , \last$104 , \ready$105 , \ready$106 , \ready$107 , pid
);
  reg \$auto$verilog_backend.cc:2083:dump_module$13  = 0;
  wire \$171 ;
  wire \$173 ;
  wire \$175 ;
  wire \$177 ;
  wire \$179 ;
  wire \$181 ;
  wire \$183 ;
  wire \$185 ;
  wire \$187 ;
  wire \$189 ;
  wire \$192 ;
  wire \$194 ;
  wire \$196 ;
  wire \$199 ;
  wire \$202 ;
  wire \$205 ;
  wire \$207 ;
  wire \$210 ;
  wire \$213 ;
  wire \$216 ;
  wire \$218 ;
  wire \$221 ;
  wire \$224 ;
  wire \$227 ;
  reg \$sample$s$valid$usb$1  = 1'h0;
  reg \$sample$s$valid$usb$1$220  = 1'h0;
  wire \$sample$s$valid$usb$1$220$next ;
  reg \$sample$s$valid$usb$1$223  = 1'h0;
  wire \$sample$s$valid$usb$1$223$next ;
  reg \$sample$s$valid$usb$1$226  = 1'h0;
  wire \$sample$s$valid$usb$1$226$next ;
  wire \$sample$s$valid$usb$1$next ;
  input ack;
  wire ack;
  output \ack$11 ;
  wire \ack$11 ;
  wire \ack$131 ;
  output \ack$3 ;
  wire \ack$3 ;
  output \ack$32 ;
  wire \ack$32 ;
  output \ack$58 ;
  wire \ack$58 ;
  input \ack$77 ;
  wire \ack$77 ;
  input \ack$78 ;
  wire \ack$78 ;
  input \ack$79 ;
  wire \ack$79 ;
  input \ack$80 ;
  wire \ack$80 ;
  input [6:0] active_address;
  wire [6:0] active_address;
  wire [6:0] \active_address$112 ;
  wire [6:0] \active_address$126 ;
  wire [6:0] \active_address$144 ;
  wire [6:0] \active_address$158 ;
  input [7:0] active_config;
  wire [7:0] active_config;
  wire [7:0] \active_config$125 ;
  wire [7:0] \active_config$143 ;
  wire [7:0] \active_config$157 ;
  output [7:0] \active_config$31 ;
  wire [7:0] \active_config$31 ;
  input [6:0] address;
  wire [6:0] address;
  wire [6:0] \address$136 ;
  output [6:0] \address$16 ;
  wire [6:0] \address$16 ;
  output [6:0] \address$37 ;
  wire [6:0] \address$37 ;
  output [6:0] \address$63 ;
  wire [6:0] \address$63 ;
  output address_changed;
  reg address_changed;
  wire \address_changed$159 ;
  wire \address_changed$160 ;
  wire \address_changed$161 ;
  input \address_changed$73 ;
  wire \address_changed$73 ;
  output config_changed;
  reg config_changed;
  wire \config_changed$165 ;
  wire \config_changed$166 ;
  wire \config_changed$167 ;
  input \config_changed$75 ;
  wire \config_changed$75 ;
  input [15:0] crc;
  wire [15:0] crc;
  wire [15:0] \crc$113 ;
  wire [15:0] \crc$127 ;
  wire [15:0] \crc$145 ;
  output [15:0] \crc$7 ;
  wire [15:0] \crc$7 ;
  input [3:0] endpoint;
  wire [3:0] endpoint;
  output [3:0] \endpoint$17 ;
  wire [3:0] \endpoint$17 ;
  output [3:0] \endpoint$38 ;
  wire [3:0] \endpoint$38 ;
  output [3:0] \endpoint$47 ;
  wire [3:0] \endpoint$47 ;
  output [3:0] \endpoint$64 ;
  wire [3:0] \endpoint$64 ;
  output first;
  wire first;
  input \first$100 ;
  wire \first$100 ;
  input \first$101 ;
  wire \first$101 ;
  input \first$99 ;
  wire \first$99 ;
  input [10:0] frame;
  wire [10:0] frame;
  wire [10:0] \frame$138 ;
  output [10:0] \frame$20 ;
  wire [10:0] \frame$20 ;
  output [10:0] \frame$41 ;
  wire [10:0] \frame$41 ;
  output [10:0] \frame$67 ;
  wire [10:0] \frame$67 ;
  input is_in;
  wire is_in;
  wire \is_in$140 ;
  output \is_in$22 ;
  wire \is_in$22 ;
  output \is_in$43 ;
  wire \is_in$43 ;
  output \is_in$69 ;
  wire \is_in$69 ;
  input is_out;
  wire is_out;
  output \is_out$23 ;
  wire \is_out$23 ;
  output \is_out$44 ;
  wire \is_out$44 ;
  output \is_out$49 ;
  wire \is_out$49 ;
  output \is_out$70 ;
  wire \is_out$70 ;
  input is_ping;
  wire is_ping;
  output \is_ping$25 ;
  wire \is_ping$25 ;
  output \is_ping$46 ;
  wire \is_ping$46 ;
  output \is_ping$50 ;
  wire \is_ping$50 ;
  output \is_ping$72 ;
  wire \is_ping$72 ;
  input is_setup;
  wire is_setup;
  wire \is_setup$141 ;
  output \is_setup$24 ;
  wire \is_setup$24 ;
  output \is_setup$45 ;
  wire \is_setup$45 ;
  output \is_setup$71 ;
  wire \is_setup$71 ;
  output last;
  wire last;
  input \last$102 ;
  wire \last$102 ;
  input \last$103 ;
  wire \last$103 ;
  input \last$104 ;
  wire \last$104 ;
  input nak;
  wire nak;
  output \nak$12 ;
  wire \nak$12 ;
  wire \nak$132 ;
  output \nak$33 ;
  wire \nak$33 ;
  output \nak$4 ;
  wire \nak$4 ;
  output \nak$59 ;
  wire \nak$59 ;
  input \nak$81 ;
  wire \nak$81 ;
  input \nak$82 ;
  wire \nak$82 ;
  input \nak$83 ;
  wire \nak$83 ;
  input \nak$84 ;
  wire \nak$84 ;
  output [6:0] new_address;
  reg [6:0] new_address;
  wire [6:0] \new_address$162 ;
  wire [6:0] \new_address$163 ;
  wire [6:0] \new_address$164 ;
  input [6:0] \new_address$74 ;
  wire [6:0] \new_address$74 ;
  output [7:0] new_config;
  reg [7:0] new_config;
  wire [7:0] \new_config$168 ;
  wire [7:0] \new_config$169 ;
  wire [7:0] \new_config$170 ;
  input [7:0] \new_config$76 ;
  wire [7:0] \new_config$76 ;
  input new_frame;
  wire new_frame;
  wire \new_frame$139 ;
  output \new_frame$21 ;
  wire \new_frame$21 ;
  output \new_frame$42 ;
  wire \new_frame$42 ;
  output \new_frame$68 ;
  wire \new_frame$68 ;
  input new_token;
  wire new_token;
  wire \new_token$137 ;
  output \new_token$18 ;
  wire \new_token$18 ;
  output \new_token$39 ;
  wire \new_token$39 ;
  output \new_token$65 ;
  wire \new_token$65 ;
  input next;
  wire next;
  wire \next$118 ;
  wire \next$150 ;
  output \next$27 ;
  wire \next$27 ;
  output \next$52 ;
  wire \next$52 ;
  input nyet;
  wire nyet;
  wire \nyet$134 ;
  output \nyet$14 ;
  wire \nyet$14 ;
  output \nyet$35 ;
  wire \nyet$35 ;
  output \nyet$61 ;
  wire \nyet$61 ;
  input [7:0] payload;
  wire [7:0] payload;
  wire [7:0] \payload$119 ;
  wire [7:0] \payload$151 ;
  output [7:0] \payload$2 ;
  wire [7:0] \payload$2 ;
  output [7:0] \payload$28 ;
  wire [7:0] \payload$28 ;
  output [7:0] \payload$53 ;
  wire [7:0] \payload$53 ;
  input [7:0] \payload$96 ;
  wire [7:0] \payload$96 ;
  input [7:0] \payload$97 ;
  wire [7:0] \payload$97 ;
  input [7:0] \payload$98 ;
  wire [7:0] \payload$98 ;
  input [3:0] pid;
  wire [3:0] pid;
  wire [3:0] \pid$135 ;
  output [3:0] \pid$15 ;
  wire [3:0] \pid$15 ;
  output [3:0] \pid$36 ;
  wire [3:0] \pid$36 ;
  output [3:0] \pid$62 ;
  wire [3:0] \pid$62 ;
  input ready;
  wire ready;
  output \ready$105 ;
  wire \ready$105 ;
  output \ready$106 ;
  wire \ready$106 ;
  output \ready$107 ;
  wire \ready$107 ;
  input ready_for_response;
  wire ready_for_response;
  output \ready_for_response$19 ;
  wire \ready_for_response$19 ;
  output \ready_for_response$40 ;
  wire \ready_for_response$40 ;
  output \ready_for_response$48 ;
  wire \ready_for_response$48 ;
  output \ready_for_response$66 ;
  wire \ready_for_response$66 ;
  input rx_complete;
  wire rx_complete;
  wire \rx_complete$109 ;
  wire \rx_complete$120 ;
  wire \rx_complete$152 ;
  output \rx_complete$54 ;
  wire \rx_complete$54 ;
  input rx_invalid;
  wire rx_invalid;
  wire \rx_invalid$110 ;
  wire \rx_invalid$122 ;
  wire \rx_invalid$154 ;
  output \rx_invalid$56 ;
  wire \rx_invalid$56 ;
  input [1:0] rx_pid_toggle;
  wire [1:0] rx_pid_toggle;
  wire [1:0] \rx_pid_toggle$111 ;
  wire [1:0] \rx_pid_toggle$123 ;
  wire [1:0] \rx_pid_toggle$155 ;
  output [1:0] \rx_pid_toggle$57 ;
  wire [1:0] \rx_pid_toggle$57 ;
  input rx_ready_for_response;
  wire rx_ready_for_response;
  wire \rx_ready_for_response$121 ;
  wire \rx_ready_for_response$153 ;
  output \rx_ready_for_response$29 ;
  wire \rx_ready_for_response$29 ;
  output \rx_ready_for_response$55 ;
  wire \rx_ready_for_response$55 ;
  input rx_timeout;
  wire rx_timeout;
  output \rx_timeout$10 ;
  wire \rx_timeout$10 ;
  wire \rx_timeout$116 ;
  wire \rx_timeout$130 ;
  wire \rx_timeout$148 ;
  input [1:0] speed;
  wire [1:0] speed;
  wire [1:0] \speed$124 ;
  wire [1:0] \speed$142 ;
  wire [1:0] \speed$156 ;
  output [1:0] \speed$30 ;
  wire [1:0] \speed$30 ;
  input stall;
  wire stall;
  output \stall$13 ;
  wire \stall$13 ;
  wire \stall$133 ;
  wire \stall$191 ;
  output \stall$34 ;
  wire \stall$34 ;
  output \stall$5 ;
  wire \stall$5 ;
  output \stall$60 ;
  wire \stall$60 ;
  input \stall$85 ;
  wire \stall$85 ;
  input \stall$86 ;
  wire \stall$86 ;
  input \stall$87 ;
  wire \stall$87 ;
  output start;
  wire start;
  wire \start$198 ;
  wire \start$201 ;
  wire \start$204 ;
  wire \start$209 ;
  wire \start$212 ;
  wire \start$215 ;
  output \start$6 ;
  wire \start$6 ;
  input \start$88 ;
  wire \start$88 ;
  input \start$89 ;
  wire \start$89 ;
  input tx_allowed;
  wire tx_allowed;
  wire \tx_allowed$114 ;
  wire \tx_allowed$128 ;
  wire \tx_allowed$146 ;
  output \tx_allowed$8 ;
  wire \tx_allowed$8 ;
  wire tx_mux_first;
  wire tx_mux_last;
  wire [7:0] tx_mux_payload;
  wire tx_mux_ready;
  wire tx_mux_valid;
  wire \tx_mux_valid$108 ;
  output [1:0] tx_pid_toggle;
  reg [1:0] tx_pid_toggle;
  wire [1:0] \tx_pid_toggle$229 ;
  input [1:0] \tx_pid_toggle$93 ;
  wire [1:0] \tx_pid_toggle$93 ;
  input [1:0] \tx_pid_toggle$94 ;
  wire [1:0] \tx_pid_toggle$94 ;
  input [1:0] \tx_pid_toggle$95 ;
  wire [1:0] \tx_pid_toggle$95 ;
  input tx_timeout;
  wire tx_timeout;
  wire \tx_timeout$115 ;
  wire \tx_timeout$129 ;
  wire \tx_timeout$147 ;
  output \tx_timeout$9 ;
  wire \tx_timeout$9 ;
  input usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  input valid;
  wire valid;
  output \valid$1 ;
  wire \valid$1 ;
  wire \valid$117 ;
  wire \valid$149 ;
  output \valid$26 ;
  wire \valid$26 ;
  output \valid$51 ;
  wire \valid$51 ;
  input \valid$90 ;
  wire \valid$90 ;
  input \valid$91 ;
  wire \valid$91 ;
  input \valid$92 ;
  wire \valid$92 ;
  assign \$173  = \$171  |  \ack$78 ;
  assign \$175  = \$173  |  \ack$79 ;
  assign \$177  = \$175  |  \ack$80 ;
  assign \$181  = \$179  |  \nak$82 ;
  assign \$183  = \$181  |  \nak$83 ;
  assign \$185  = \$183  |  \nak$84 ;
  assign \$189  = \$187  |  \stall$86 ;
  assign \$194  = \$192  |  \stall$87 ;
  assign \$218  = \valid$90  |  \$sample$s$valid$usb$1 ;
  assign \$221  = \valid$91  |  \$sample$s$valid$usb$1$220 ;
  assign \$227  = \valid$92  |  \$sample$s$valid$usb$1$226 ;
  always @(posedge usb_clk)
    \$sample$s$valid$usb$1  <= \$sample$s$valid$usb$1$next ;
  always @(posedge usb_clk)
    \$sample$s$valid$usb$1$220  <= \$sample$s$valid$usb$1$220$next ;
  always @(posedge usb_clk)
    \$sample$s$valid$usb$1$223  <= 1'h0;
  always @(posedge usb_clk)
    \$sample$s$valid$usb$1$226  <= \$sample$s$valid$usb$1$226$next ;
  tx_mux tx_mux (
    .first(tx_mux_first),
    .\first$10 (\first$101 ),
    .\first$8 (\first$99 ),
    .\first$9 (\first$100 ),
    .last(tx_mux_last),
    .\last$11 (\last$102 ),
    .\last$12 (\last$103 ),
    .\last$13 (\last$104 ),
    .payload(tx_mux_payload),
    .\payload$5 (\payload$96 ),
    .\payload$6 (\payload$97 ),
    .\payload$7 (\payload$98 ),
    .ready(tx_mux_ready),
    .\ready$14 (\ready$105 ),
    .\ready$15 (\ready$106 ),
    .\ready$16 (\ready$107 ),
    .valid(tx_mux_valid),
    .\valid$1 (\valid$90 ),
    .\valid$2 (\valid$91 ),
    .\valid$3 (1'h0),
    .\valid$4 (\valid$92 )
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$13 ) begin end
    address_changed = 1'h0;
    casez ({ \address_changed$161 , \address_changed$160 , \address_changed$159 , \address_changed$73  })
      4'b???1:
          address_changed = \address_changed$73 ;
      4'b??1?:
          address_changed = 1'h0;
      4'b?1??:
          address_changed = 1'h0;
      4'b1???:
          address_changed = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$13 ) begin end
    new_address = 7'h00;
    casez ({ \address_changed$161 , \address_changed$160 , \address_changed$159 , \address_changed$73  })
      4'b???1:
          new_address = \new_address$74 ;
      4'b??1?:
          new_address = 7'h00;
      4'b?1??:
          new_address = 7'h00;
      4'b1???:
          new_address = 7'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$13 ) begin end
    config_changed = 1'h0;
    casez ({ \config_changed$167 , \config_changed$166 , \config_changed$165 , \config_changed$75  })
      4'b???1:
          config_changed = \config_changed$75 ;
      4'b??1?:
          config_changed = 1'h0;
      4'b?1??:
          config_changed = 1'h0;
      4'b1???:
          config_changed = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$13 ) begin end
    new_config = 8'h00;
    casez ({ \config_changed$167 , \config_changed$166 , \config_changed$165 , \config_changed$75  })
      4'b???1:
          new_config = \new_config$76 ;
      4'b??1?:
          new_config = 8'h00;
      4'b?1??:
          new_config = 8'h00;
      4'b1???:
          new_config = 8'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$13 ) begin end
    tx_pid_toggle = 2'h0;
    casez ({ \$227 , \$224 , \$221 , \$218  })
      4'b???1:
          tx_pid_toggle = \tx_pid_toggle$93 ;
      4'b??1?:
          tx_pid_toggle = \tx_pid_toggle$94 ;
      4'b?1??:
          tx_pid_toggle = 2'h0;
      4'b1???:
          tx_pid_toggle = \tx_pid_toggle$95 ;
    endcase
  end
  assign \tx_mux_valid$108  = 1'h0;
  assign \address_changed$159  = 1'h0;
  assign \address_changed$160  = 1'h0;
  assign \address_changed$161  = 1'h0;
  assign \new_address$162  = 7'h00;
  assign \new_address$163  = 7'h00;
  assign \new_address$164  = 7'h00;
  assign \config_changed$165  = 1'h0;
  assign \config_changed$166  = 1'h0;
  assign \config_changed$167  = 1'h0;
  assign \new_config$168  = 8'h00;
  assign \new_config$169  = 8'h00;
  assign \new_config$170  = 8'h00;
  assign \stall$191  = 1'h0;
  assign \start$198  = 1'h0;
  assign \start$201  = 1'h0;
  assign \start$204  = 1'h0;
  assign \start$209  = 1'h0;
  assign \start$212  = 1'h0;
  assign \start$215  = 1'h0;
  assign \tx_pid_toggle$229  = 2'h0;
  assign \$sample$s$valid$usb$1$226$next  = \valid$92 ;
  assign \$sample$s$valid$usb$1$223$next  = 1'h0;
  assign \$sample$s$valid$usb$1$220$next  = \valid$91 ;
  assign \$sample$s$valid$usb$1$next  = \valid$90 ;
  assign \start$6  = \$216 ;
  assign start = \$205 ;
  assign \stall$5  = \$194 ;
  assign \nak$4  = \$185 ;
  assign \ack$3  = \$177 ;
  assign tx_mux_ready = ready;
  assign \payload$2  = tx_mux_payload;
  assign last = tx_mux_last;
  assign first = tx_mux_first;
  assign \valid$1  = tx_mux_valid;
  assign \active_address$158  = active_address;
  assign \active_config$157  = active_config;
  assign \speed$156  = speed;
  assign \rx_pid_toggle$155  = rx_pid_toggle;
  assign \rx_invalid$154  = rx_invalid;
  assign \rx_ready_for_response$153  = rx_ready_for_response;
  assign \rx_complete$152  = rx_complete;
  assign \payload$151  = payload;
  assign \next$150  = next;
  assign \valid$149  = valid;
  assign \is_ping$72  = is_ping;
  assign \is_setup$71  = is_setup;
  assign \is_out$70  = is_out;
  assign \is_in$69  = is_in;
  assign \new_frame$68  = new_frame;
  assign \frame$67  = frame;
  assign \ready_for_response$66  = ready_for_response;
  assign \new_token$65  = new_token;
  assign \endpoint$64  = endpoint;
  assign \address$63  = address;
  assign \pid$62  = pid;
  assign \nyet$61  = nyet;
  assign \stall$60  = stall;
  assign \nak$59  = nak;
  assign \ack$58  = ack;
  assign \rx_timeout$148  = rx_timeout;
  assign \tx_timeout$147  = tx_timeout;
  assign \tx_allowed$146  = tx_allowed;
  assign \crc$145  = crc;
  assign \active_address$144  = active_address;
  assign \active_config$143  = active_config;
  assign \speed$142  = speed;
  assign \rx_pid_toggle$57  = rx_pid_toggle;
  assign \rx_invalid$56  = rx_invalid;
  assign \rx_ready_for_response$55  = rx_ready_for_response;
  assign \rx_complete$54  = rx_complete;
  assign \payload$53  = payload;
  assign \next$52  = next;
  assign \valid$51  = valid;
  assign \is_ping$50  = is_ping;
  assign \is_setup$141  = is_setup;
  assign \is_out$49  = is_out;
  assign \is_in$140  = is_in;
  assign \new_frame$139  = new_frame;
  assign \frame$138  = frame;
  assign \ready_for_response$48  = ready_for_response;
  assign \new_token$137  = new_token;
  assign \endpoint$47  = endpoint;
  assign \address$136  = address;
  assign \pid$135  = pid;
  assign \nyet$134  = nyet;
  assign \stall$133  = stall;
  assign \nak$132  = nak;
  assign \ack$131  = ack;
  assign \rx_timeout$130  = rx_timeout;
  assign \tx_timeout$129  = tx_timeout;
  assign \tx_allowed$128  = tx_allowed;
  assign \crc$127  = crc;
  assign \active_address$126  = active_address;
  assign \active_config$125  = active_config;
  assign \speed$124  = speed;
  assign \rx_pid_toggle$123  = rx_pid_toggle;
  assign \rx_invalid$122  = rx_invalid;
  assign \rx_ready_for_response$121  = rx_ready_for_response;
  assign \rx_complete$120  = rx_complete;
  assign \payload$119  = payload;
  assign \next$118  = next;
  assign \valid$117  = valid;
  assign \is_ping$46  = is_ping;
  assign \is_setup$45  = is_setup;
  assign \is_out$44  = is_out;
  assign \is_in$43  = is_in;
  assign \new_frame$42  = new_frame;
  assign \frame$41  = frame;
  assign \ready_for_response$40  = ready_for_response;
  assign \new_token$39  = new_token;
  assign \endpoint$38  = endpoint;
  assign \address$37  = address;
  assign \pid$36  = pid;
  assign \nyet$35  = nyet;
  assign \stall$34  = stall;
  assign \nak$33  = nak;
  assign \ack$32  = ack;
  assign \rx_timeout$116  = rx_timeout;
  assign \tx_timeout$115  = tx_timeout;
  assign \tx_allowed$114  = tx_allowed;
  assign \crc$113  = crc;
  assign \active_address$112  = active_address;
  assign \active_config$31  = active_config;
  assign \speed$30  = speed;
  assign \rx_pid_toggle$111  = rx_pid_toggle;
  assign \rx_invalid$110  = rx_invalid;
  assign \rx_ready_for_response$29  = rx_ready_for_response;
  assign \rx_complete$109  = rx_complete;
  assign \payload$28  = payload;
  assign \next$27  = next;
  assign \valid$26  = valid;
  assign \is_ping$25  = is_ping;
  assign \is_setup$24  = is_setup;
  assign \is_out$23  = is_out;
  assign \is_in$22  = is_in;
  assign \new_frame$21  = new_frame;
  assign \frame$20  = frame;
  assign \ready_for_response$19  = ready_for_response;
  assign \new_token$18  = new_token;
  assign \endpoint$17  = endpoint;
  assign \address$16  = address;
  assign \pid$15  = pid;
  assign \nyet$14  = nyet;
  assign \stall$13  = stall;
  assign \nak$12  = nak;
  assign \ack$11  = ack;
  assign \rx_timeout$10  = rx_timeout;
  assign \tx_timeout$9  = tx_timeout;
  assign \tx_allowed$8  = tx_allowed;
  assign \crc$7  = crc;
  assign \$171  = \ack$77 ;
  assign \$179  = \nak$81 ;
  assign \$187  = \stall$85 ;
  assign \$192  = \$189 ;
  assign \$196  = \start$88 ;
  assign \$199  = \start$88 ;
  assign \$202  = \start$88 ;
  assign \$205  = \start$88 ;
  assign \$207  = \start$89 ;
  assign \$210  = \start$89 ;
  assign \$213  = \start$89 ;
  assign \$216  = \start$89 ;
  assign \$224  = \$sample$s$valid$usb$1$223 ;
endmodule
module fifo(usb_clk, write_data, write_en, full, write_commit, write_discard, space_available, empty, read_data, read_en, read_commit, usb_rst);
  reg \$auto$verilog_backend.cc:2083:dump_module$14  = 0;
  wire \$11 ;
  wire \$13 ;
  wire \$15 ;
  wire [10:0] \$17 ;
  wire [10:0] \$18 ;
  wire \$2 ;
  wire \$20 ;
  wire \$22 ;
  wire \$24 ;
  wire \$26 ;
  wire \$28 ;
  wire \$30 ;
  wire [11:0] \$32 ;
  wire [10:0] \$33 ;
  wire [11:0] \$35 ;
  wire [11:0] \$37 ;
  wire [10:0] \$38 ;
  wire \$4 ;
  wire [11:0] \$40 ;
  wire \$42 ;
  wire \$6 ;
  wire [10:0] \$8 ;
  wire [10:0] \$9 ;
  reg [9:0] committed_read_pointer = 10'h000;
  reg [9:0] \committed_read_pointer$next ;
  reg [9:0] committed_write_pointer = 10'h000;
  reg [9:0] \committed_write_pointer$next ;
  reg [9:0] current_read_pointer = 10'h000;
  reg [9:0] \current_read_pointer$next ;
  reg [9:0] current_write_pointer = 10'h000;
  reg [9:0] \current_write_pointer$next ;
  output empty;
  wire empty;
  output full;
  wire full;
  reg [9:0] next_read_pointer;
  reg [9:0] next_write_pointer;
  input read_commit;
  wire read_commit;
  output [9:0] read_data;
  wire [9:0] read_data;
  wire read_discard;
  input read_en;
  wire read_en;
  reg [9:0] rx_fifo_r_addr;
  wire [9:0] rx_fifo_r_data;
  wire [9:0] rx_fifo_w_addr;
  wire [9:0] rx_fifo_w_data;
  wire rx_fifo_w_en;
  output [9:0] space_available;
  reg [9:0] space_available;
  input usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  input write_commit;
  wire write_commit;
  input [9:0] write_data;
  wire [9:0] write_data;
  input write_discard;
  wire write_discard;
  input write_en;
  wire write_en;
  reg [9:0] rx_fifo [1023:0];
  initial begin
    rx_fifo[0] = 10'h000;
    rx_fifo[1] = 10'h000;
    rx_fifo[2] = 10'h000;
    rx_fifo[3] = 10'h000;
    rx_fifo[4] = 10'h000;
    rx_fifo[5] = 10'h000;
    rx_fifo[6] = 10'h000;
    rx_fifo[7] = 10'h000;
    rx_fifo[8] = 10'h000;
    rx_fifo[9] = 10'h000;
    rx_fifo[10] = 10'h000;
    rx_fifo[11] = 10'h000;
    rx_fifo[12] = 10'h000;
    rx_fifo[13] = 10'h000;
    rx_fifo[14] = 10'h000;
    rx_fifo[15] = 10'h000;
    rx_fifo[16] = 10'h000;
    rx_fifo[17] = 10'h000;
    rx_fifo[18] = 10'h000;
    rx_fifo[19] = 10'h000;
    rx_fifo[20] = 10'h000;
    rx_fifo[21] = 10'h000;
    rx_fifo[22] = 10'h000;
    rx_fifo[23] = 10'h000;
    rx_fifo[24] = 10'h000;
    rx_fifo[25] = 10'h000;
    rx_fifo[26] = 10'h000;
    rx_fifo[27] = 10'h000;
    rx_fifo[28] = 10'h000;
    rx_fifo[29] = 10'h000;
    rx_fifo[30] = 10'h000;
    rx_fifo[31] = 10'h000;
    rx_fifo[32] = 10'h000;
    rx_fifo[33] = 10'h000;
    rx_fifo[34] = 10'h000;
    rx_fifo[35] = 10'h000;
    rx_fifo[36] = 10'h000;
    rx_fifo[37] = 10'h000;
    rx_fifo[38] = 10'h000;
    rx_fifo[39] = 10'h000;
    rx_fifo[40] = 10'h000;
    rx_fifo[41] = 10'h000;
    rx_fifo[42] = 10'h000;
    rx_fifo[43] = 10'h000;
    rx_fifo[44] = 10'h000;
    rx_fifo[45] = 10'h000;
    rx_fifo[46] = 10'h000;
    rx_fifo[47] = 10'h000;
    rx_fifo[48] = 10'h000;
    rx_fifo[49] = 10'h000;
    rx_fifo[50] = 10'h000;
    rx_fifo[51] = 10'h000;
    rx_fifo[52] = 10'h000;
    rx_fifo[53] = 10'h000;
    rx_fifo[54] = 10'h000;
    rx_fifo[55] = 10'h000;
    rx_fifo[56] = 10'h000;
    rx_fifo[57] = 10'h000;
    rx_fifo[58] = 10'h000;
    rx_fifo[59] = 10'h000;
    rx_fifo[60] = 10'h000;
    rx_fifo[61] = 10'h000;
    rx_fifo[62] = 10'h000;
    rx_fifo[63] = 10'h000;
    rx_fifo[64] = 10'h000;
    rx_fifo[65] = 10'h000;
    rx_fifo[66] = 10'h000;
    rx_fifo[67] = 10'h000;
    rx_fifo[68] = 10'h000;
    rx_fifo[69] = 10'h000;
    rx_fifo[70] = 10'h000;
    rx_fifo[71] = 10'h000;
    rx_fifo[72] = 10'h000;
    rx_fifo[73] = 10'h000;
    rx_fifo[74] = 10'h000;
    rx_fifo[75] = 10'h000;
    rx_fifo[76] = 10'h000;
    rx_fifo[77] = 10'h000;
    rx_fifo[78] = 10'h000;
    rx_fifo[79] = 10'h000;
    rx_fifo[80] = 10'h000;
    rx_fifo[81] = 10'h000;
    rx_fifo[82] = 10'h000;
    rx_fifo[83] = 10'h000;
    rx_fifo[84] = 10'h000;
    rx_fifo[85] = 10'h000;
    rx_fifo[86] = 10'h000;
    rx_fifo[87] = 10'h000;
    rx_fifo[88] = 10'h000;
    rx_fifo[89] = 10'h000;
    rx_fifo[90] = 10'h000;
    rx_fifo[91] = 10'h000;
    rx_fifo[92] = 10'h000;
    rx_fifo[93] = 10'h000;
    rx_fifo[94] = 10'h000;
    rx_fifo[95] = 10'h000;
    rx_fifo[96] = 10'h000;
    rx_fifo[97] = 10'h000;
    rx_fifo[98] = 10'h000;
    rx_fifo[99] = 10'h000;
    rx_fifo[100] = 10'h000;
    rx_fifo[101] = 10'h000;
    rx_fifo[102] = 10'h000;
    rx_fifo[103] = 10'h000;
    rx_fifo[104] = 10'h000;
    rx_fifo[105] = 10'h000;
    rx_fifo[106] = 10'h000;
    rx_fifo[107] = 10'h000;
    rx_fifo[108] = 10'h000;
    rx_fifo[109] = 10'h000;
    rx_fifo[110] = 10'h000;
    rx_fifo[111] = 10'h000;
    rx_fifo[112] = 10'h000;
    rx_fifo[113] = 10'h000;
    rx_fifo[114] = 10'h000;
    rx_fifo[115] = 10'h000;
    rx_fifo[116] = 10'h000;
    rx_fifo[117] = 10'h000;
    rx_fifo[118] = 10'h000;
    rx_fifo[119] = 10'h000;
    rx_fifo[120] = 10'h000;
    rx_fifo[121] = 10'h000;
    rx_fifo[122] = 10'h000;
    rx_fifo[123] = 10'h000;
    rx_fifo[124] = 10'h000;
    rx_fifo[125] = 10'h000;
    rx_fifo[126] = 10'h000;
    rx_fifo[127] = 10'h000;
    rx_fifo[128] = 10'h000;
    rx_fifo[129] = 10'h000;
    rx_fifo[130] = 10'h000;
    rx_fifo[131] = 10'h000;
    rx_fifo[132] = 10'h000;
    rx_fifo[133] = 10'h000;
    rx_fifo[134] = 10'h000;
    rx_fifo[135] = 10'h000;
    rx_fifo[136] = 10'h000;
    rx_fifo[137] = 10'h000;
    rx_fifo[138] = 10'h000;
    rx_fifo[139] = 10'h000;
    rx_fifo[140] = 10'h000;
    rx_fifo[141] = 10'h000;
    rx_fifo[142] = 10'h000;
    rx_fifo[143] = 10'h000;
    rx_fifo[144] = 10'h000;
    rx_fifo[145] = 10'h000;
    rx_fifo[146] = 10'h000;
    rx_fifo[147] = 10'h000;
    rx_fifo[148] = 10'h000;
    rx_fifo[149] = 10'h000;
    rx_fifo[150] = 10'h000;
    rx_fifo[151] = 10'h000;
    rx_fifo[152] = 10'h000;
    rx_fifo[153] = 10'h000;
    rx_fifo[154] = 10'h000;
    rx_fifo[155] = 10'h000;
    rx_fifo[156] = 10'h000;
    rx_fifo[157] = 10'h000;
    rx_fifo[158] = 10'h000;
    rx_fifo[159] = 10'h000;
    rx_fifo[160] = 10'h000;
    rx_fifo[161] = 10'h000;
    rx_fifo[162] = 10'h000;
    rx_fifo[163] = 10'h000;
    rx_fifo[164] = 10'h000;
    rx_fifo[165] = 10'h000;
    rx_fifo[166] = 10'h000;
    rx_fifo[167] = 10'h000;
    rx_fifo[168] = 10'h000;
    rx_fifo[169] = 10'h000;
    rx_fifo[170] = 10'h000;
    rx_fifo[171] = 10'h000;
    rx_fifo[172] = 10'h000;
    rx_fifo[173] = 10'h000;
    rx_fifo[174] = 10'h000;
    rx_fifo[175] = 10'h000;
    rx_fifo[176] = 10'h000;
    rx_fifo[177] = 10'h000;
    rx_fifo[178] = 10'h000;
    rx_fifo[179] = 10'h000;
    rx_fifo[180] = 10'h000;
    rx_fifo[181] = 10'h000;
    rx_fifo[182] = 10'h000;
    rx_fifo[183] = 10'h000;
    rx_fifo[184] = 10'h000;
    rx_fifo[185] = 10'h000;
    rx_fifo[186] = 10'h000;
    rx_fifo[187] = 10'h000;
    rx_fifo[188] = 10'h000;
    rx_fifo[189] = 10'h000;
    rx_fifo[190] = 10'h000;
    rx_fifo[191] = 10'h000;
    rx_fifo[192] = 10'h000;
    rx_fifo[193] = 10'h000;
    rx_fifo[194] = 10'h000;
    rx_fifo[195] = 10'h000;
    rx_fifo[196] = 10'h000;
    rx_fifo[197] = 10'h000;
    rx_fifo[198] = 10'h000;
    rx_fifo[199] = 10'h000;
    rx_fifo[200] = 10'h000;
    rx_fifo[201] = 10'h000;
    rx_fifo[202] = 10'h000;
    rx_fifo[203] = 10'h000;
    rx_fifo[204] = 10'h000;
    rx_fifo[205] = 10'h000;
    rx_fifo[206] = 10'h000;
    rx_fifo[207] = 10'h000;
    rx_fifo[208] = 10'h000;
    rx_fifo[209] = 10'h000;
    rx_fifo[210] = 10'h000;
    rx_fifo[211] = 10'h000;
    rx_fifo[212] = 10'h000;
    rx_fifo[213] = 10'h000;
    rx_fifo[214] = 10'h000;
    rx_fifo[215] = 10'h000;
    rx_fifo[216] = 10'h000;
    rx_fifo[217] = 10'h000;
    rx_fifo[218] = 10'h000;
    rx_fifo[219] = 10'h000;
    rx_fifo[220] = 10'h000;
    rx_fifo[221] = 10'h000;
    rx_fifo[222] = 10'h000;
    rx_fifo[223] = 10'h000;
    rx_fifo[224] = 10'h000;
    rx_fifo[225] = 10'h000;
    rx_fifo[226] = 10'h000;
    rx_fifo[227] = 10'h000;
    rx_fifo[228] = 10'h000;
    rx_fifo[229] = 10'h000;
    rx_fifo[230] = 10'h000;
    rx_fifo[231] = 10'h000;
    rx_fifo[232] = 10'h000;
    rx_fifo[233] = 10'h000;
    rx_fifo[234] = 10'h000;
    rx_fifo[235] = 10'h000;
    rx_fifo[236] = 10'h000;
    rx_fifo[237] = 10'h000;
    rx_fifo[238] = 10'h000;
    rx_fifo[239] = 10'h000;
    rx_fifo[240] = 10'h000;
    rx_fifo[241] = 10'h000;
    rx_fifo[242] = 10'h000;
    rx_fifo[243] = 10'h000;
    rx_fifo[244] = 10'h000;
    rx_fifo[245] = 10'h000;
    rx_fifo[246] = 10'h000;
    rx_fifo[247] = 10'h000;
    rx_fifo[248] = 10'h000;
    rx_fifo[249] = 10'h000;
    rx_fifo[250] = 10'h000;
    rx_fifo[251] = 10'h000;
    rx_fifo[252] = 10'h000;
    rx_fifo[253] = 10'h000;
    rx_fifo[254] = 10'h000;
    rx_fifo[255] = 10'h000;
    rx_fifo[256] = 10'h000;
    rx_fifo[257] = 10'h000;
    rx_fifo[258] = 10'h000;
    rx_fifo[259] = 10'h000;
    rx_fifo[260] = 10'h000;
    rx_fifo[261] = 10'h000;
    rx_fifo[262] = 10'h000;
    rx_fifo[263] = 10'h000;
    rx_fifo[264] = 10'h000;
    rx_fifo[265] = 10'h000;
    rx_fifo[266] = 10'h000;
    rx_fifo[267] = 10'h000;
    rx_fifo[268] = 10'h000;
    rx_fifo[269] = 10'h000;
    rx_fifo[270] = 10'h000;
    rx_fifo[271] = 10'h000;
    rx_fifo[272] = 10'h000;
    rx_fifo[273] = 10'h000;
    rx_fifo[274] = 10'h000;
    rx_fifo[275] = 10'h000;
    rx_fifo[276] = 10'h000;
    rx_fifo[277] = 10'h000;
    rx_fifo[278] = 10'h000;
    rx_fifo[279] = 10'h000;
    rx_fifo[280] = 10'h000;
    rx_fifo[281] = 10'h000;
    rx_fifo[282] = 10'h000;
    rx_fifo[283] = 10'h000;
    rx_fifo[284] = 10'h000;
    rx_fifo[285] = 10'h000;
    rx_fifo[286] = 10'h000;
    rx_fifo[287] = 10'h000;
    rx_fifo[288] = 10'h000;
    rx_fifo[289] = 10'h000;
    rx_fifo[290] = 10'h000;
    rx_fifo[291] = 10'h000;
    rx_fifo[292] = 10'h000;
    rx_fifo[293] = 10'h000;
    rx_fifo[294] = 10'h000;
    rx_fifo[295] = 10'h000;
    rx_fifo[296] = 10'h000;
    rx_fifo[297] = 10'h000;
    rx_fifo[298] = 10'h000;
    rx_fifo[299] = 10'h000;
    rx_fifo[300] = 10'h000;
    rx_fifo[301] = 10'h000;
    rx_fifo[302] = 10'h000;
    rx_fifo[303] = 10'h000;
    rx_fifo[304] = 10'h000;
    rx_fifo[305] = 10'h000;
    rx_fifo[306] = 10'h000;
    rx_fifo[307] = 10'h000;
    rx_fifo[308] = 10'h000;
    rx_fifo[309] = 10'h000;
    rx_fifo[310] = 10'h000;
    rx_fifo[311] = 10'h000;
    rx_fifo[312] = 10'h000;
    rx_fifo[313] = 10'h000;
    rx_fifo[314] = 10'h000;
    rx_fifo[315] = 10'h000;
    rx_fifo[316] = 10'h000;
    rx_fifo[317] = 10'h000;
    rx_fifo[318] = 10'h000;
    rx_fifo[319] = 10'h000;
    rx_fifo[320] = 10'h000;
    rx_fifo[321] = 10'h000;
    rx_fifo[322] = 10'h000;
    rx_fifo[323] = 10'h000;
    rx_fifo[324] = 10'h000;
    rx_fifo[325] = 10'h000;
    rx_fifo[326] = 10'h000;
    rx_fifo[327] = 10'h000;
    rx_fifo[328] = 10'h000;
    rx_fifo[329] = 10'h000;
    rx_fifo[330] = 10'h000;
    rx_fifo[331] = 10'h000;
    rx_fifo[332] = 10'h000;
    rx_fifo[333] = 10'h000;
    rx_fifo[334] = 10'h000;
    rx_fifo[335] = 10'h000;
    rx_fifo[336] = 10'h000;
    rx_fifo[337] = 10'h000;
    rx_fifo[338] = 10'h000;
    rx_fifo[339] = 10'h000;
    rx_fifo[340] = 10'h000;
    rx_fifo[341] = 10'h000;
    rx_fifo[342] = 10'h000;
    rx_fifo[343] = 10'h000;
    rx_fifo[344] = 10'h000;
    rx_fifo[345] = 10'h000;
    rx_fifo[346] = 10'h000;
    rx_fifo[347] = 10'h000;
    rx_fifo[348] = 10'h000;
    rx_fifo[349] = 10'h000;
    rx_fifo[350] = 10'h000;
    rx_fifo[351] = 10'h000;
    rx_fifo[352] = 10'h000;
    rx_fifo[353] = 10'h000;
    rx_fifo[354] = 10'h000;
    rx_fifo[355] = 10'h000;
    rx_fifo[356] = 10'h000;
    rx_fifo[357] = 10'h000;
    rx_fifo[358] = 10'h000;
    rx_fifo[359] = 10'h000;
    rx_fifo[360] = 10'h000;
    rx_fifo[361] = 10'h000;
    rx_fifo[362] = 10'h000;
    rx_fifo[363] = 10'h000;
    rx_fifo[364] = 10'h000;
    rx_fifo[365] = 10'h000;
    rx_fifo[366] = 10'h000;
    rx_fifo[367] = 10'h000;
    rx_fifo[368] = 10'h000;
    rx_fifo[369] = 10'h000;
    rx_fifo[370] = 10'h000;
    rx_fifo[371] = 10'h000;
    rx_fifo[372] = 10'h000;
    rx_fifo[373] = 10'h000;
    rx_fifo[374] = 10'h000;
    rx_fifo[375] = 10'h000;
    rx_fifo[376] = 10'h000;
    rx_fifo[377] = 10'h000;
    rx_fifo[378] = 10'h000;
    rx_fifo[379] = 10'h000;
    rx_fifo[380] = 10'h000;
    rx_fifo[381] = 10'h000;
    rx_fifo[382] = 10'h000;
    rx_fifo[383] = 10'h000;
    rx_fifo[384] = 10'h000;
    rx_fifo[385] = 10'h000;
    rx_fifo[386] = 10'h000;
    rx_fifo[387] = 10'h000;
    rx_fifo[388] = 10'h000;
    rx_fifo[389] = 10'h000;
    rx_fifo[390] = 10'h000;
    rx_fifo[391] = 10'h000;
    rx_fifo[392] = 10'h000;
    rx_fifo[393] = 10'h000;
    rx_fifo[394] = 10'h000;
    rx_fifo[395] = 10'h000;
    rx_fifo[396] = 10'h000;
    rx_fifo[397] = 10'h000;
    rx_fifo[398] = 10'h000;
    rx_fifo[399] = 10'h000;
    rx_fifo[400] = 10'h000;
    rx_fifo[401] = 10'h000;
    rx_fifo[402] = 10'h000;
    rx_fifo[403] = 10'h000;
    rx_fifo[404] = 10'h000;
    rx_fifo[405] = 10'h000;
    rx_fifo[406] = 10'h000;
    rx_fifo[407] = 10'h000;
    rx_fifo[408] = 10'h000;
    rx_fifo[409] = 10'h000;
    rx_fifo[410] = 10'h000;
    rx_fifo[411] = 10'h000;
    rx_fifo[412] = 10'h000;
    rx_fifo[413] = 10'h000;
    rx_fifo[414] = 10'h000;
    rx_fifo[415] = 10'h000;
    rx_fifo[416] = 10'h000;
    rx_fifo[417] = 10'h000;
    rx_fifo[418] = 10'h000;
    rx_fifo[419] = 10'h000;
    rx_fifo[420] = 10'h000;
    rx_fifo[421] = 10'h000;
    rx_fifo[422] = 10'h000;
    rx_fifo[423] = 10'h000;
    rx_fifo[424] = 10'h000;
    rx_fifo[425] = 10'h000;
    rx_fifo[426] = 10'h000;
    rx_fifo[427] = 10'h000;
    rx_fifo[428] = 10'h000;
    rx_fifo[429] = 10'h000;
    rx_fifo[430] = 10'h000;
    rx_fifo[431] = 10'h000;
    rx_fifo[432] = 10'h000;
    rx_fifo[433] = 10'h000;
    rx_fifo[434] = 10'h000;
    rx_fifo[435] = 10'h000;
    rx_fifo[436] = 10'h000;
    rx_fifo[437] = 10'h000;
    rx_fifo[438] = 10'h000;
    rx_fifo[439] = 10'h000;
    rx_fifo[440] = 10'h000;
    rx_fifo[441] = 10'h000;
    rx_fifo[442] = 10'h000;
    rx_fifo[443] = 10'h000;
    rx_fifo[444] = 10'h000;
    rx_fifo[445] = 10'h000;
    rx_fifo[446] = 10'h000;
    rx_fifo[447] = 10'h000;
    rx_fifo[448] = 10'h000;
    rx_fifo[449] = 10'h000;
    rx_fifo[450] = 10'h000;
    rx_fifo[451] = 10'h000;
    rx_fifo[452] = 10'h000;
    rx_fifo[453] = 10'h000;
    rx_fifo[454] = 10'h000;
    rx_fifo[455] = 10'h000;
    rx_fifo[456] = 10'h000;
    rx_fifo[457] = 10'h000;
    rx_fifo[458] = 10'h000;
    rx_fifo[459] = 10'h000;
    rx_fifo[460] = 10'h000;
    rx_fifo[461] = 10'h000;
    rx_fifo[462] = 10'h000;
    rx_fifo[463] = 10'h000;
    rx_fifo[464] = 10'h000;
    rx_fifo[465] = 10'h000;
    rx_fifo[466] = 10'h000;
    rx_fifo[467] = 10'h000;
    rx_fifo[468] = 10'h000;
    rx_fifo[469] = 10'h000;
    rx_fifo[470] = 10'h000;
    rx_fifo[471] = 10'h000;
    rx_fifo[472] = 10'h000;
    rx_fifo[473] = 10'h000;
    rx_fifo[474] = 10'h000;
    rx_fifo[475] = 10'h000;
    rx_fifo[476] = 10'h000;
    rx_fifo[477] = 10'h000;
    rx_fifo[478] = 10'h000;
    rx_fifo[479] = 10'h000;
    rx_fifo[480] = 10'h000;
    rx_fifo[481] = 10'h000;
    rx_fifo[482] = 10'h000;
    rx_fifo[483] = 10'h000;
    rx_fifo[484] = 10'h000;
    rx_fifo[485] = 10'h000;
    rx_fifo[486] = 10'h000;
    rx_fifo[487] = 10'h000;
    rx_fifo[488] = 10'h000;
    rx_fifo[489] = 10'h000;
    rx_fifo[490] = 10'h000;
    rx_fifo[491] = 10'h000;
    rx_fifo[492] = 10'h000;
    rx_fifo[493] = 10'h000;
    rx_fifo[494] = 10'h000;
    rx_fifo[495] = 10'h000;
    rx_fifo[496] = 10'h000;
    rx_fifo[497] = 10'h000;
    rx_fifo[498] = 10'h000;
    rx_fifo[499] = 10'h000;
    rx_fifo[500] = 10'h000;
    rx_fifo[501] = 10'h000;
    rx_fifo[502] = 10'h000;
    rx_fifo[503] = 10'h000;
    rx_fifo[504] = 10'h000;
    rx_fifo[505] = 10'h000;
    rx_fifo[506] = 10'h000;
    rx_fifo[507] = 10'h000;
    rx_fifo[508] = 10'h000;
    rx_fifo[509] = 10'h000;
    rx_fifo[510] = 10'h000;
    rx_fifo[511] = 10'h000;
    rx_fifo[512] = 10'h000;
    rx_fifo[513] = 10'h000;
    rx_fifo[514] = 10'h000;
    rx_fifo[515] = 10'h000;
    rx_fifo[516] = 10'h000;
    rx_fifo[517] = 10'h000;
    rx_fifo[518] = 10'h000;
    rx_fifo[519] = 10'h000;
    rx_fifo[520] = 10'h000;
    rx_fifo[521] = 10'h000;
    rx_fifo[522] = 10'h000;
    rx_fifo[523] = 10'h000;
    rx_fifo[524] = 10'h000;
    rx_fifo[525] = 10'h000;
    rx_fifo[526] = 10'h000;
    rx_fifo[527] = 10'h000;
    rx_fifo[528] = 10'h000;
    rx_fifo[529] = 10'h000;
    rx_fifo[530] = 10'h000;
    rx_fifo[531] = 10'h000;
    rx_fifo[532] = 10'h000;
    rx_fifo[533] = 10'h000;
    rx_fifo[534] = 10'h000;
    rx_fifo[535] = 10'h000;
    rx_fifo[536] = 10'h000;
    rx_fifo[537] = 10'h000;
    rx_fifo[538] = 10'h000;
    rx_fifo[539] = 10'h000;
    rx_fifo[540] = 10'h000;
    rx_fifo[541] = 10'h000;
    rx_fifo[542] = 10'h000;
    rx_fifo[543] = 10'h000;
    rx_fifo[544] = 10'h000;
    rx_fifo[545] = 10'h000;
    rx_fifo[546] = 10'h000;
    rx_fifo[547] = 10'h000;
    rx_fifo[548] = 10'h000;
    rx_fifo[549] = 10'h000;
    rx_fifo[550] = 10'h000;
    rx_fifo[551] = 10'h000;
    rx_fifo[552] = 10'h000;
    rx_fifo[553] = 10'h000;
    rx_fifo[554] = 10'h000;
    rx_fifo[555] = 10'h000;
    rx_fifo[556] = 10'h000;
    rx_fifo[557] = 10'h000;
    rx_fifo[558] = 10'h000;
    rx_fifo[559] = 10'h000;
    rx_fifo[560] = 10'h000;
    rx_fifo[561] = 10'h000;
    rx_fifo[562] = 10'h000;
    rx_fifo[563] = 10'h000;
    rx_fifo[564] = 10'h000;
    rx_fifo[565] = 10'h000;
    rx_fifo[566] = 10'h000;
    rx_fifo[567] = 10'h000;
    rx_fifo[568] = 10'h000;
    rx_fifo[569] = 10'h000;
    rx_fifo[570] = 10'h000;
    rx_fifo[571] = 10'h000;
    rx_fifo[572] = 10'h000;
    rx_fifo[573] = 10'h000;
    rx_fifo[574] = 10'h000;
    rx_fifo[575] = 10'h000;
    rx_fifo[576] = 10'h000;
    rx_fifo[577] = 10'h000;
    rx_fifo[578] = 10'h000;
    rx_fifo[579] = 10'h000;
    rx_fifo[580] = 10'h000;
    rx_fifo[581] = 10'h000;
    rx_fifo[582] = 10'h000;
    rx_fifo[583] = 10'h000;
    rx_fifo[584] = 10'h000;
    rx_fifo[585] = 10'h000;
    rx_fifo[586] = 10'h000;
    rx_fifo[587] = 10'h000;
    rx_fifo[588] = 10'h000;
    rx_fifo[589] = 10'h000;
    rx_fifo[590] = 10'h000;
    rx_fifo[591] = 10'h000;
    rx_fifo[592] = 10'h000;
    rx_fifo[593] = 10'h000;
    rx_fifo[594] = 10'h000;
    rx_fifo[595] = 10'h000;
    rx_fifo[596] = 10'h000;
    rx_fifo[597] = 10'h000;
    rx_fifo[598] = 10'h000;
    rx_fifo[599] = 10'h000;
    rx_fifo[600] = 10'h000;
    rx_fifo[601] = 10'h000;
    rx_fifo[602] = 10'h000;
    rx_fifo[603] = 10'h000;
    rx_fifo[604] = 10'h000;
    rx_fifo[605] = 10'h000;
    rx_fifo[606] = 10'h000;
    rx_fifo[607] = 10'h000;
    rx_fifo[608] = 10'h000;
    rx_fifo[609] = 10'h000;
    rx_fifo[610] = 10'h000;
    rx_fifo[611] = 10'h000;
    rx_fifo[612] = 10'h000;
    rx_fifo[613] = 10'h000;
    rx_fifo[614] = 10'h000;
    rx_fifo[615] = 10'h000;
    rx_fifo[616] = 10'h000;
    rx_fifo[617] = 10'h000;
    rx_fifo[618] = 10'h000;
    rx_fifo[619] = 10'h000;
    rx_fifo[620] = 10'h000;
    rx_fifo[621] = 10'h000;
    rx_fifo[622] = 10'h000;
    rx_fifo[623] = 10'h000;
    rx_fifo[624] = 10'h000;
    rx_fifo[625] = 10'h000;
    rx_fifo[626] = 10'h000;
    rx_fifo[627] = 10'h000;
    rx_fifo[628] = 10'h000;
    rx_fifo[629] = 10'h000;
    rx_fifo[630] = 10'h000;
    rx_fifo[631] = 10'h000;
    rx_fifo[632] = 10'h000;
    rx_fifo[633] = 10'h000;
    rx_fifo[634] = 10'h000;
    rx_fifo[635] = 10'h000;
    rx_fifo[636] = 10'h000;
    rx_fifo[637] = 10'h000;
    rx_fifo[638] = 10'h000;
    rx_fifo[639] = 10'h000;
    rx_fifo[640] = 10'h000;
    rx_fifo[641] = 10'h000;
    rx_fifo[642] = 10'h000;
    rx_fifo[643] = 10'h000;
    rx_fifo[644] = 10'h000;
    rx_fifo[645] = 10'h000;
    rx_fifo[646] = 10'h000;
    rx_fifo[647] = 10'h000;
    rx_fifo[648] = 10'h000;
    rx_fifo[649] = 10'h000;
    rx_fifo[650] = 10'h000;
    rx_fifo[651] = 10'h000;
    rx_fifo[652] = 10'h000;
    rx_fifo[653] = 10'h000;
    rx_fifo[654] = 10'h000;
    rx_fifo[655] = 10'h000;
    rx_fifo[656] = 10'h000;
    rx_fifo[657] = 10'h000;
    rx_fifo[658] = 10'h000;
    rx_fifo[659] = 10'h000;
    rx_fifo[660] = 10'h000;
    rx_fifo[661] = 10'h000;
    rx_fifo[662] = 10'h000;
    rx_fifo[663] = 10'h000;
    rx_fifo[664] = 10'h000;
    rx_fifo[665] = 10'h000;
    rx_fifo[666] = 10'h000;
    rx_fifo[667] = 10'h000;
    rx_fifo[668] = 10'h000;
    rx_fifo[669] = 10'h000;
    rx_fifo[670] = 10'h000;
    rx_fifo[671] = 10'h000;
    rx_fifo[672] = 10'h000;
    rx_fifo[673] = 10'h000;
    rx_fifo[674] = 10'h000;
    rx_fifo[675] = 10'h000;
    rx_fifo[676] = 10'h000;
    rx_fifo[677] = 10'h000;
    rx_fifo[678] = 10'h000;
    rx_fifo[679] = 10'h000;
    rx_fifo[680] = 10'h000;
    rx_fifo[681] = 10'h000;
    rx_fifo[682] = 10'h000;
    rx_fifo[683] = 10'h000;
    rx_fifo[684] = 10'h000;
    rx_fifo[685] = 10'h000;
    rx_fifo[686] = 10'h000;
    rx_fifo[687] = 10'h000;
    rx_fifo[688] = 10'h000;
    rx_fifo[689] = 10'h000;
    rx_fifo[690] = 10'h000;
    rx_fifo[691] = 10'h000;
    rx_fifo[692] = 10'h000;
    rx_fifo[693] = 10'h000;
    rx_fifo[694] = 10'h000;
    rx_fifo[695] = 10'h000;
    rx_fifo[696] = 10'h000;
    rx_fifo[697] = 10'h000;
    rx_fifo[698] = 10'h000;
    rx_fifo[699] = 10'h000;
    rx_fifo[700] = 10'h000;
    rx_fifo[701] = 10'h000;
    rx_fifo[702] = 10'h000;
    rx_fifo[703] = 10'h000;
    rx_fifo[704] = 10'h000;
    rx_fifo[705] = 10'h000;
    rx_fifo[706] = 10'h000;
    rx_fifo[707] = 10'h000;
    rx_fifo[708] = 10'h000;
    rx_fifo[709] = 10'h000;
    rx_fifo[710] = 10'h000;
    rx_fifo[711] = 10'h000;
    rx_fifo[712] = 10'h000;
    rx_fifo[713] = 10'h000;
    rx_fifo[714] = 10'h000;
    rx_fifo[715] = 10'h000;
    rx_fifo[716] = 10'h000;
    rx_fifo[717] = 10'h000;
    rx_fifo[718] = 10'h000;
    rx_fifo[719] = 10'h000;
    rx_fifo[720] = 10'h000;
    rx_fifo[721] = 10'h000;
    rx_fifo[722] = 10'h000;
    rx_fifo[723] = 10'h000;
    rx_fifo[724] = 10'h000;
    rx_fifo[725] = 10'h000;
    rx_fifo[726] = 10'h000;
    rx_fifo[727] = 10'h000;
    rx_fifo[728] = 10'h000;
    rx_fifo[729] = 10'h000;
    rx_fifo[730] = 10'h000;
    rx_fifo[731] = 10'h000;
    rx_fifo[732] = 10'h000;
    rx_fifo[733] = 10'h000;
    rx_fifo[734] = 10'h000;
    rx_fifo[735] = 10'h000;
    rx_fifo[736] = 10'h000;
    rx_fifo[737] = 10'h000;
    rx_fifo[738] = 10'h000;
    rx_fifo[739] = 10'h000;
    rx_fifo[740] = 10'h000;
    rx_fifo[741] = 10'h000;
    rx_fifo[742] = 10'h000;
    rx_fifo[743] = 10'h000;
    rx_fifo[744] = 10'h000;
    rx_fifo[745] = 10'h000;
    rx_fifo[746] = 10'h000;
    rx_fifo[747] = 10'h000;
    rx_fifo[748] = 10'h000;
    rx_fifo[749] = 10'h000;
    rx_fifo[750] = 10'h000;
    rx_fifo[751] = 10'h000;
    rx_fifo[752] = 10'h000;
    rx_fifo[753] = 10'h000;
    rx_fifo[754] = 10'h000;
    rx_fifo[755] = 10'h000;
    rx_fifo[756] = 10'h000;
    rx_fifo[757] = 10'h000;
    rx_fifo[758] = 10'h000;
    rx_fifo[759] = 10'h000;
    rx_fifo[760] = 10'h000;
    rx_fifo[761] = 10'h000;
    rx_fifo[762] = 10'h000;
    rx_fifo[763] = 10'h000;
    rx_fifo[764] = 10'h000;
    rx_fifo[765] = 10'h000;
    rx_fifo[766] = 10'h000;
    rx_fifo[767] = 10'h000;
    rx_fifo[768] = 10'h000;
    rx_fifo[769] = 10'h000;
    rx_fifo[770] = 10'h000;
    rx_fifo[771] = 10'h000;
    rx_fifo[772] = 10'h000;
    rx_fifo[773] = 10'h000;
    rx_fifo[774] = 10'h000;
    rx_fifo[775] = 10'h000;
    rx_fifo[776] = 10'h000;
    rx_fifo[777] = 10'h000;
    rx_fifo[778] = 10'h000;
    rx_fifo[779] = 10'h000;
    rx_fifo[780] = 10'h000;
    rx_fifo[781] = 10'h000;
    rx_fifo[782] = 10'h000;
    rx_fifo[783] = 10'h000;
    rx_fifo[784] = 10'h000;
    rx_fifo[785] = 10'h000;
    rx_fifo[786] = 10'h000;
    rx_fifo[787] = 10'h000;
    rx_fifo[788] = 10'h000;
    rx_fifo[789] = 10'h000;
    rx_fifo[790] = 10'h000;
    rx_fifo[791] = 10'h000;
    rx_fifo[792] = 10'h000;
    rx_fifo[793] = 10'h000;
    rx_fifo[794] = 10'h000;
    rx_fifo[795] = 10'h000;
    rx_fifo[796] = 10'h000;
    rx_fifo[797] = 10'h000;
    rx_fifo[798] = 10'h000;
    rx_fifo[799] = 10'h000;
    rx_fifo[800] = 10'h000;
    rx_fifo[801] = 10'h000;
    rx_fifo[802] = 10'h000;
    rx_fifo[803] = 10'h000;
    rx_fifo[804] = 10'h000;
    rx_fifo[805] = 10'h000;
    rx_fifo[806] = 10'h000;
    rx_fifo[807] = 10'h000;
    rx_fifo[808] = 10'h000;
    rx_fifo[809] = 10'h000;
    rx_fifo[810] = 10'h000;
    rx_fifo[811] = 10'h000;
    rx_fifo[812] = 10'h000;
    rx_fifo[813] = 10'h000;
    rx_fifo[814] = 10'h000;
    rx_fifo[815] = 10'h000;
    rx_fifo[816] = 10'h000;
    rx_fifo[817] = 10'h000;
    rx_fifo[818] = 10'h000;
    rx_fifo[819] = 10'h000;
    rx_fifo[820] = 10'h000;
    rx_fifo[821] = 10'h000;
    rx_fifo[822] = 10'h000;
    rx_fifo[823] = 10'h000;
    rx_fifo[824] = 10'h000;
    rx_fifo[825] = 10'h000;
    rx_fifo[826] = 10'h000;
    rx_fifo[827] = 10'h000;
    rx_fifo[828] = 10'h000;
    rx_fifo[829] = 10'h000;
    rx_fifo[830] = 10'h000;
    rx_fifo[831] = 10'h000;
    rx_fifo[832] = 10'h000;
    rx_fifo[833] = 10'h000;
    rx_fifo[834] = 10'h000;
    rx_fifo[835] = 10'h000;
    rx_fifo[836] = 10'h000;
    rx_fifo[837] = 10'h000;
    rx_fifo[838] = 10'h000;
    rx_fifo[839] = 10'h000;
    rx_fifo[840] = 10'h000;
    rx_fifo[841] = 10'h000;
    rx_fifo[842] = 10'h000;
    rx_fifo[843] = 10'h000;
    rx_fifo[844] = 10'h000;
    rx_fifo[845] = 10'h000;
    rx_fifo[846] = 10'h000;
    rx_fifo[847] = 10'h000;
    rx_fifo[848] = 10'h000;
    rx_fifo[849] = 10'h000;
    rx_fifo[850] = 10'h000;
    rx_fifo[851] = 10'h000;
    rx_fifo[852] = 10'h000;
    rx_fifo[853] = 10'h000;
    rx_fifo[854] = 10'h000;
    rx_fifo[855] = 10'h000;
    rx_fifo[856] = 10'h000;
    rx_fifo[857] = 10'h000;
    rx_fifo[858] = 10'h000;
    rx_fifo[859] = 10'h000;
    rx_fifo[860] = 10'h000;
    rx_fifo[861] = 10'h000;
    rx_fifo[862] = 10'h000;
    rx_fifo[863] = 10'h000;
    rx_fifo[864] = 10'h000;
    rx_fifo[865] = 10'h000;
    rx_fifo[866] = 10'h000;
    rx_fifo[867] = 10'h000;
    rx_fifo[868] = 10'h000;
    rx_fifo[869] = 10'h000;
    rx_fifo[870] = 10'h000;
    rx_fifo[871] = 10'h000;
    rx_fifo[872] = 10'h000;
    rx_fifo[873] = 10'h000;
    rx_fifo[874] = 10'h000;
    rx_fifo[875] = 10'h000;
    rx_fifo[876] = 10'h000;
    rx_fifo[877] = 10'h000;
    rx_fifo[878] = 10'h000;
    rx_fifo[879] = 10'h000;
    rx_fifo[880] = 10'h000;
    rx_fifo[881] = 10'h000;
    rx_fifo[882] = 10'h000;
    rx_fifo[883] = 10'h000;
    rx_fifo[884] = 10'h000;
    rx_fifo[885] = 10'h000;
    rx_fifo[886] = 10'h000;
    rx_fifo[887] = 10'h000;
    rx_fifo[888] = 10'h000;
    rx_fifo[889] = 10'h000;
    rx_fifo[890] = 10'h000;
    rx_fifo[891] = 10'h000;
    rx_fifo[892] = 10'h000;
    rx_fifo[893] = 10'h000;
    rx_fifo[894] = 10'h000;
    rx_fifo[895] = 10'h000;
    rx_fifo[896] = 10'h000;
    rx_fifo[897] = 10'h000;
    rx_fifo[898] = 10'h000;
    rx_fifo[899] = 10'h000;
    rx_fifo[900] = 10'h000;
    rx_fifo[901] = 10'h000;
    rx_fifo[902] = 10'h000;
    rx_fifo[903] = 10'h000;
    rx_fifo[904] = 10'h000;
    rx_fifo[905] = 10'h000;
    rx_fifo[906] = 10'h000;
    rx_fifo[907] = 10'h000;
    rx_fifo[908] = 10'h000;
    rx_fifo[909] = 10'h000;
    rx_fifo[910] = 10'h000;
    rx_fifo[911] = 10'h000;
    rx_fifo[912] = 10'h000;
    rx_fifo[913] = 10'h000;
    rx_fifo[914] = 10'h000;
    rx_fifo[915] = 10'h000;
    rx_fifo[916] = 10'h000;
    rx_fifo[917] = 10'h000;
    rx_fifo[918] = 10'h000;
    rx_fifo[919] = 10'h000;
    rx_fifo[920] = 10'h000;
    rx_fifo[921] = 10'h000;
    rx_fifo[922] = 10'h000;
    rx_fifo[923] = 10'h000;
    rx_fifo[924] = 10'h000;
    rx_fifo[925] = 10'h000;
    rx_fifo[926] = 10'h000;
    rx_fifo[927] = 10'h000;
    rx_fifo[928] = 10'h000;
    rx_fifo[929] = 10'h000;
    rx_fifo[930] = 10'h000;
    rx_fifo[931] = 10'h000;
    rx_fifo[932] = 10'h000;
    rx_fifo[933] = 10'h000;
    rx_fifo[934] = 10'h000;
    rx_fifo[935] = 10'h000;
    rx_fifo[936] = 10'h000;
    rx_fifo[937] = 10'h000;
    rx_fifo[938] = 10'h000;
    rx_fifo[939] = 10'h000;
    rx_fifo[940] = 10'h000;
    rx_fifo[941] = 10'h000;
    rx_fifo[942] = 10'h000;
    rx_fifo[943] = 10'h000;
    rx_fifo[944] = 10'h000;
    rx_fifo[945] = 10'h000;
    rx_fifo[946] = 10'h000;
    rx_fifo[947] = 10'h000;
    rx_fifo[948] = 10'h000;
    rx_fifo[949] = 10'h000;
    rx_fifo[950] = 10'h000;
    rx_fifo[951] = 10'h000;
    rx_fifo[952] = 10'h000;
    rx_fifo[953] = 10'h000;
    rx_fifo[954] = 10'h000;
    rx_fifo[955] = 10'h000;
    rx_fifo[956] = 10'h000;
    rx_fifo[957] = 10'h000;
    rx_fifo[958] = 10'h000;
    rx_fifo[959] = 10'h000;
    rx_fifo[960] = 10'h000;
    rx_fifo[961] = 10'h000;
    rx_fifo[962] = 10'h000;
    rx_fifo[963] = 10'h000;
    rx_fifo[964] = 10'h000;
    rx_fifo[965] = 10'h000;
    rx_fifo[966] = 10'h000;
    rx_fifo[967] = 10'h000;
    rx_fifo[968] = 10'h000;
    rx_fifo[969] = 10'h000;
    rx_fifo[970] = 10'h000;
    rx_fifo[971] = 10'h000;
    rx_fifo[972] = 10'h000;
    rx_fifo[973] = 10'h000;
    rx_fifo[974] = 10'h000;
    rx_fifo[975] = 10'h000;
    rx_fifo[976] = 10'h000;
    rx_fifo[977] = 10'h000;
    rx_fifo[978] = 10'h000;
    rx_fifo[979] = 10'h000;
    rx_fifo[980] = 10'h000;
    rx_fifo[981] = 10'h000;
    rx_fifo[982] = 10'h000;
    rx_fifo[983] = 10'h000;
    rx_fifo[984] = 10'h000;
    rx_fifo[985] = 10'h000;
    rx_fifo[986] = 10'h000;
    rx_fifo[987] = 10'h000;
    rx_fifo[988] = 10'h000;
    rx_fifo[989] = 10'h000;
    rx_fifo[990] = 10'h000;
    rx_fifo[991] = 10'h000;
    rx_fifo[992] = 10'h000;
    rx_fifo[993] = 10'h000;
    rx_fifo[994] = 10'h000;
    rx_fifo[995] = 10'h000;
    rx_fifo[996] = 10'h000;
    rx_fifo[997] = 10'h000;
    rx_fifo[998] = 10'h000;
    rx_fifo[999] = 10'h000;
    rx_fifo[1000] = 10'h000;
    rx_fifo[1001] = 10'h000;
    rx_fifo[1002] = 10'h000;
    rx_fifo[1003] = 10'h000;
    rx_fifo[1004] = 10'h000;
    rx_fifo[1005] = 10'h000;
    rx_fifo[1006] = 10'h000;
    rx_fifo[1007] = 10'h000;
    rx_fifo[1008] = 10'h000;
    rx_fifo[1009] = 10'h000;
    rx_fifo[1010] = 10'h000;
    rx_fifo[1011] = 10'h000;
    rx_fifo[1012] = 10'h000;
    rx_fifo[1013] = 10'h000;
    rx_fifo[1014] = 10'h000;
    rx_fifo[1015] = 10'h000;
    rx_fifo[1016] = 10'h000;
    rx_fifo[1017] = 10'h000;
    rx_fifo[1018] = 10'h000;
    rx_fifo[1019] = 10'h000;
    rx_fifo[1020] = 10'h000;
    rx_fifo[1021] = 10'h000;
    rx_fifo[1022] = 10'h000;
    rx_fifo[1023] = 10'h000;
  end
  always @(posedge usb_clk) begin
    if (rx_fifo_w_en)
      rx_fifo[rx_fifo_w_addr] <= rx_fifo_w_data;
  end
  reg [9:0] _0_;
  always @(posedge usb_clk) begin
    _0_ <= rx_fifo_r_addr;
  end
  assign rx_fifo_r_data = rx_fifo[_0_];
  assign \$9  = current_write_pointer +  1'h1;
  assign \$11  = ~  full;
  assign \$13  = write_en &  \$11 ;
  assign \$15  = current_read_pointer ==  10'h3ff;
  assign \$18  = current_read_pointer +  1'h1;
  assign \$20  = ~  empty;
  assign \$22  = read_en &  \$20 ;
  assign \$24  = ~  empty;
  assign \$26  = read_en &  \$24 ;
  assign \$28  = current_read_pointer ==  committed_write_pointer;
  assign \$2  = ~  full;
  assign \$30  = committed_read_pointer <=  current_write_pointer;
  assign \$33  = current_write_pointer -  committed_read_pointer;
  assign \$35  = 10'h3ff -  \$33 ;
  assign \$38  = committed_read_pointer -  current_write_pointer;
  assign \$40  = \$38  -  1'h1;
  assign \$42  = next_write_pointer ==  committed_read_pointer;
  always @(posedge usb_clk)
    current_write_pointer <= \current_write_pointer$next ;
  always @(posedge usb_clk)
    committed_write_pointer <= \committed_write_pointer$next ;
  always @(posedge usb_clk)
    current_read_pointer <= \current_read_pointer$next ;
  always @(posedge usb_clk)
    committed_read_pointer <= \committed_read_pointer$next ;
  assign \$4  = write_en &  \$2 ;
  assign \$6  = current_write_pointer ==  10'h3ff;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$14 ) begin end
    \committed_read_pointer$next  = committed_read_pointer;
    casez (read_commit)
      1'h1:
          \committed_read_pointer$next  = current_read_pointer;
    endcase
    casez (usb_rst)
      1'h1:
          \committed_read_pointer$next  = 10'h000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$14 ) begin end
    casez ({ \$30 , full })
      2'b?1:
          space_available = 10'h000;
      2'b1?:
          space_available = \$35 [9:0];
      default:
          space_available = \$40 [9:0];
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$14 ) begin end
    casez (\$6 )
      1'h1:
          next_write_pointer = 10'h000;
      default:
          next_write_pointer = \$9 [9:0];
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$14 ) begin end
    \current_write_pointer$next  = current_write_pointer;
    casez (\$13 )
      1'h1:
          \current_write_pointer$next  = next_write_pointer;
    endcase
    casez (write_discard)
      1'h1:
          \current_write_pointer$next  = committed_write_pointer;
    endcase
    casez (usb_rst)
      1'h1:
          \current_write_pointer$next  = 10'h000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$14 ) begin end
    \committed_write_pointer$next  = committed_write_pointer;
    casez (write_commit)
      1'h1:
          \committed_write_pointer$next  = current_write_pointer;
    endcase
    casez (usb_rst)
      1'h1:
          \committed_write_pointer$next  = 10'h000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$14 ) begin end
    casez (\$15 )
      1'h1:
          next_read_pointer = 10'h000;
      default:
          next_read_pointer = \$18 [9:0];
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$14 ) begin end
    casez (\$22 )
      1'h1:
          rx_fifo_r_addr = next_read_pointer;
      default:
          rx_fifo_r_addr = current_read_pointer;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$14 ) begin end
    \current_read_pointer$next  = current_read_pointer;
    casez (\$26 )
      1'h1:
          \current_read_pointer$next  = next_read_pointer;
    endcase
    casez (read_discard)
      1'h1:
          \current_read_pointer$next  = committed_read_pointer;
    endcase
    casez (usb_rst)
      1'h1:
          \current_read_pointer$next  = 10'h000;
    endcase
  end
  assign \$8  = \$9 ;
  assign \$17  = \$18 ;
  assign \$32  = \$35 ;
  assign \$37  = \$40 ;
  assign read_discard = 1'h0;
  assign full = \$42 ;
  assign empty = \$28 ;
  assign rx_fifo_w_addr = current_write_pointer;
  assign rx_fifo_w_en = \$4 ;
  assign rx_fifo_w_data = write_data;
  assign read_data = rx_fifo_r_data;
endmodule
module get_descriptor(usb_clk, value, length, start_position, valid, first, last, payload, ready, stall, start, usb_rst);
  reg \$auto$verilog_backend.cc:2083:dump_module$15  = 0;
  wire \$10 ;
  wire [16:0] \$100 ;
  wire \$102 ;
  wire \$104 ;
  wire \$107 ;
  wire [16:0] \$108 ;
  wire [16:0] \$11 ;
  wire \$110 ;
  wire [16:0] \$112 ;
  wire \$114 ;
  wire \$116 ;
  wire [7:0] \$119 ;
  wire [2:0] \$120 ;
  wire [6:0] \$122 ;
  wire \$125 ;
  wire [16:0] \$127 ;
  wire \$129 ;
  wire \$13 ;
  wire [16:0] \$131 ;
  wire \$133 ;
  wire \$135 ;
  wire [16:0] \$15 ;
  wire \$17 ;
  wire \$19 ;
  wire [16:0] \$22 ;
  wire [16:0] \$23 ;
  wire \$25 ;
  wire [8:0] \$27 ;
  wire [8:0] \$28 ;
  wire [16:0] \$3 ;
  wire [32:0] \$30 ;
  wire [32:0] \$31 ;
  wire [32:0] \$33 ;
  wire [6:0] \$35 ;
  wire [5:0] \$36 ;
  wire [6:0] \$38 ;
  wire \$40 ;
  wire [16:0] \$41 ;
  wire \$43 ;
  wire [16:0] \$45 ;
  wire \$47 ;
  wire \$49 ;
  wire \$5 ;
  wire [6:0] \$52 ;
  wire [6:0] \$53 ;
  wire [6:0] \$54 ;
  wire [6:0] \$56 ;
  wire \$58 ;
  wire \$60 ;
  wire \$62 ;
  wire \$64 ;
  wire [16:0] \$65 ;
  wire \$67 ;
  wire [16:0] \$69 ;
  wire [16:0] \$7 ;
  wire \$71 ;
  wire \$73 ;
  wire \$76 ;
  wire [16:0] \$77 ;
  wire \$79 ;
  wire [16:0] \$8 ;
  wire [16:0] \$81 ;
  wire \$83 ;
  wire \$85 ;
  wire [6:0] \$88 ;
  wire [6:0] \$89 ;
  wire \$91 ;
  wire \$93 ;
  wire \$95 ;
  wire [16:0] \$96 ;
  wire \$98 ;
  reg [15:0] bytes_sent = 16'h0000;
  reg [15:0] \bytes_sent$next ;
  reg [5:0] descriptor_data_base_address = 6'h00;
  reg [5:0] \descriptor_data_base_address$next ;
  reg [15:0] descriptor_length = 16'h0000;
  reg [15:0] \descriptor_length$next ;
  output first;
  reg first;
  reg [2:0] fsm_state = 3'h0;
  reg [2:0] \fsm_state$next ;
  wire [7:0] index;
  output last;
  reg last;
  input [15:0] length;
  wire [15:0] length;
  reg [15:0] \length$2  = 16'h0000;
  reg [15:0] \length$2$next ;
  output [7:0] payload;
  reg [7:0] payload;
  reg [5:0] position_in_stream = 6'h00;
  reg [5:0] \position_in_stream$next ;
  input ready;
  wire ready;
  reg [5:0] rom_r_addr;
  wire [31:0] rom_r_data;
  wire rom_r_en;
  output stall;
  reg stall;
  input start;
  wire start;
  input [10:0] start_position;
  wire [10:0] start_position;
  wire [7:0] type_number;
  input usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  output valid;
  reg valid;
  input [15:0] value;
  wire [15:0] value;
  reg [31:0] rom [57:0];
  initial begin
    rom[0] = 32'd0;
    rom[1] = 32'd65552;
    rom[2] = 32'd65556;
    rom[3] = 32'd262168;
    rom[4] = 32'd1179688;
    rom[5] = 32'd4128828;
    rom[6] = 32'd262268;
    rom[7] = 32'd917632;
    rom[8] = 32'd3932304;
    rom[9] = 32'd1835212;
    rom[10] = 32'd302055426;
    rom[11] = 32'd33554496;
    rom[12] = 32'd2671050768;
    rom[13] = 32'd258;
    rom[14] = 32'd50397184;
    rom[15] = 32'd151142144;
    rom[16] = 32'd33620096;
    rom[17] = 32'd4194894848;
    rom[18] = 32'd66050;
    rom[19] = 32'd16778532;
    rom[20] = 32'd1048837;
    rom[21] = 32'd604372993;
    rom[22] = 32'd86245632;
    rom[23] = 32'd17237379;
    rom[24] = 32'd50332171;
    rom[25] = 32'd151257344;
    rom[26] = 32'd34209792;
    rom[27] = 32'd460164;
    rom[28] = 32'd33555199;
    rom[29] = 32'd117769218;
    rom[30] = 32'd196352;
    rom[31] = 32'd67307780;
    rom[32] = 32'd235098880;
    rom[33] = 32'd1761636352;
    rom[34] = 32'd1694524672;
    rom[35] = 32'd1677721600;
    rom[36] = 32'd1006851072;
    rom[37] = 32'd1627418112;
    rom[38] = 32'd1728061440;
    rom[39] = 32'd1342206464;
    rom[40] = 32'd1761635584;
    rom[41] = 32'd1694528000;
    rom[42] = 32'd536883712;
    rom[43] = 32'd805325568;
    rom[44] = 32'd536892672;
    rom[45] = 32'd1392525824;
    rom[46] = 32'd755004416;
    rom[47] = 32'd1862282496;
    rom[48] = 32'd1929405696;
    rom[49] = 32'd1912629504;
    rom[50] = 32'd1627417600;
    rom[51] = 32'd469971200;
    rom[52] = 32'd822096896;
    rom[53] = 32'd889204992;
    rom[54] = 32'd872427776;
    rom[55] = 32'd956313856;
    rom[56] = 32'd956315648;
    rom[57] = 32'd822095872;
  end
  reg [31:0] _0_;
  always @(posedge usb_clk) begin
    _0_ <= rom[rom_r_addr];
  end
  assign rom_r_data = _0_;
  assign \$100  = bytes_sent +  1'h1;
  assign \$102  = \$100  >=  \length$2 ;
  assign \$104  = \$98  |  \$102 ;
  assign \$95  = ~  \$104 ;
  assign \$108  = descriptor_length -  1'h1;
  assign \$110  = position_in_stream ==  \$108 ;
  assign \$112  = bytes_sent +  1'h1;
  assign \$114  = \$112  >=  \length$2 ;
  assign \$116  = \$110  |  \$114 ;
  assign \$107  = ~  \$116 ;
  assign \$11  = descriptor_length -  1'h1;
  assign \$120  = 2'h3 -  position_in_stream[1:0];
  assign \$122  = \$120  *  4'h8;
  assign \$119  = rom_r_data >> \$122 ;
  assign \$125  = position_in_stream ==  start_position;
  assign \$127  = descriptor_length -  1'h1;
  assign \$129  = position_in_stream ==  \$127 ;
  assign \$131  = bytes_sent +  1'h1;
  assign \$133  = \$131  >=  \length$2 ;
  assign \$135  = \$129  |  \$133 ;
  always @(posedge usb_clk)
    \length$2  <= \length$2$next ;
  always @(posedge usb_clk)
    bytes_sent <= \bytes_sent$next ;
  always @(posedge usb_clk)
    fsm_state <= \fsm_state$next ;
  assign \$13  = position_in_stream ==  \$11 ;
  always @(posedge usb_clk)
    position_in_stream <= \position_in_stream$next ;
  always @(posedge usb_clk)
    descriptor_data_base_address <= \descriptor_data_base_address$next ;
  always @(posedge usb_clk)
    descriptor_length <= \descriptor_length$next ;
  assign \$15  = bytes_sent +  1'h1;
  assign \$17  = \$15  >=  \length$2 ;
  assign \$19  = \$13  |  \$17 ;
  assign \$10  = ~  \$19 ;
  assign \$23  = bytes_sent +  1'h1;
  assign \$25  = index >=  rom_r_data[31:16];
  assign \$28  = rom_r_data[7:2] +  index;
  assign \$31  = rom_r_data +  position_in_stream;
  assign \$38  = descriptor_data_base_address +  \$36 ;
  assign \$3  = length -  start_position;
  assign \$41  = descriptor_length -  1'h1;
  assign \$43  = position_in_stream ==  \$41 ;
  assign \$45  = bytes_sent +  1'h1;
  assign \$47  = \$45  >=  \length$2 ;
  assign \$49  = \$43  |  \$47 ;
  assign \$40  = ~  \$49 ;
  assign \$54  = position_in_stream +  1'h1;
  assign \$56  = descriptor_data_base_address +  \$53 [5:2];
  assign \$58  = type_number <=  2'h3;
  assign \$5  = \$3  <=  7'h40;
  assign \$60  = index >=  rom_r_data[31:16];
  assign \$62  = !  \length$2 ;
  assign \$65  = descriptor_length -  1'h1;
  assign \$67  = position_in_stream ==  \$65 ;
  assign \$69  = bytes_sent +  1'h1;
  assign \$71  = \$69  >=  \length$2 ;
  assign \$73  = \$67  |  \$71 ;
  assign \$64  = ~  \$73 ;
  assign \$77  = descriptor_length -  1'h1;
  assign \$79  = position_in_stream ==  \$77 ;
  assign \$81  = bytes_sent +  1'h1;
  assign \$83  = \$81  >=  \length$2 ;
  assign \$85  = \$79  |  \$83 ;
  assign \$76  = ~  \$85 ;
  assign \$8  = length -  start_position;
  assign \$89  = position_in_stream +  1'h1;
  assign \$91  = type_number <=  2'h3;
  assign \$93  = index >=  rom_r_data[31:16];
  assign \$96  = descriptor_length -  1'h1;
  assign \$98  = position_in_stream ==  \$96 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$15 ) begin end
    valid = 1'h0;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          ;
      3'h4:
          ;
      3'h5:
          valid = 1'h1;
      3'h3:
          valid = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$15 ) begin end
    payload = 8'h00;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          ;
      3'h4:
          ;
      3'h5:
          payload = \$119 ;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$15 ) begin end
    first = 1'h0;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          ;
      3'h4:
          ;
      3'h5:
          first = \$125 ;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$15 ) begin end
    last = 1'h0;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          ;
      3'h4:
          ;
      3'h5:
          last = \$135 ;
      3'h3:
          last = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$15 ) begin end
    casez (\$5 )
      1'h1:
          \length$2$next  = \$8 [15:0];
      default:
          \length$2$next  = 16'h0040;
    endcase
    casez (usb_rst)
      1'h1:
          \length$2$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$15 ) begin end
    \bytes_sent$next  = bytes_sent;
    casez (fsm_state)
      3'h0:
          \bytes_sent$next  = 16'h0000;
      3'h1:
          ;
      3'h2:
          ;
      3'h4:
          ;
      3'h5:
          casez (ready)
            1'h1:
                casez (\$10 )
                  1'h1:
                      \bytes_sent$next  = \$23 [15:0];
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \bytes_sent$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$15 ) begin end
    rom_r_addr = 6'h00;
    casez (fsm_state)
      3'h0:
          rom_r_addr = type_number[5:0];
      3'h1:
          rom_r_addr = type_number[5:0];
      3'h2:
          casez (\$25 )
            1'h1:
                ;
            default:
                rom_r_addr = \$28 [5:0];
          endcase
      3'h4:
          rom_r_addr = \$33 [5:0];
      3'h5:
        begin
          rom_r_addr = \$38 [5:0];
          casez (ready)
            1'h1:
                casez (\$40 )
                  1'h1:
                      rom_r_addr = \$56 [5:0];
                endcase
          endcase
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$15 ) begin end
    \fsm_state$next  = fsm_state;
    casez (fsm_state)
      3'h0:
          casez (start)
            1'h1:
                \fsm_state$next  = 3'h1;
          endcase
      3'h1:
          casez (\$58 )
            1'h1:
                \fsm_state$next  = 3'h2;
            default:
                \fsm_state$next  = 3'h0;
          endcase
      3'h2:
          casez (\$60 )
            1'h1:
                \fsm_state$next  = 3'h0;
            default:
                casez (\$62 )
                  1'h1:
                      \fsm_state$next  = 3'h3;
                  default:
                      \fsm_state$next  = 3'h4;
                endcase
          endcase
      3'h4:
          \fsm_state$next  = 3'h5;
      3'h5:
          casez (ready)
            1'h1:
                casez (\$64 )
                  1'h1:
                      ;
                  default:
                      \fsm_state$next  = 3'h0;
                endcase
          endcase
      3'h3:
          \fsm_state$next  = 3'h0;
    endcase
    casez (usb_rst)
      1'h1:
          \fsm_state$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$15 ) begin end
    \position_in_stream$next  = position_in_stream;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          \position_in_stream$next  = start_position[5:0];
      3'h2:
          ;
      3'h4:
          ;
      3'h5:
          casez (ready)
            1'h1:
                casez (\$76 )
                  1'h1:
                      \position_in_stream$next  = \$89 [5:0];
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \position_in_stream$next  = 6'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$15 ) begin end
    stall = 1'h0;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          casez (\$91 )
            1'h1:
                ;
            default:
                stall = 1'h1;
          endcase
      3'h2:
          casez (\$93 )
            1'h1:
                stall = 1'h1;
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$15 ) begin end
    \descriptor_data_base_address$next  = descriptor_data_base_address;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          ;
      3'h4:
          \descriptor_data_base_address$next  = rom_r_data[7:2];
      3'h5:
          casez (ready)
            1'h1:
                casez (\$95 )
                  1'h1:
                      ;
                  default:
                      \descriptor_data_base_address$next  = 6'h00;
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \descriptor_data_base_address$next  = 6'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$15 ) begin end
    \descriptor_length$next  = descriptor_length;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          ;
      3'h4:
          \descriptor_length$next  = rom_r_data[31:16];
      3'h5:
          casez (ready)
            1'h1:
                casez (\$107 )
                  1'h1:
                      ;
                  default:
                      \descriptor_length$next  = 16'h0000;
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \descriptor_length$next  = 16'h0000;
    endcase
  end
  assign \$7  = \$8 ;
  assign \$22  = \$23 ;
  assign \$27  = \$28 ;
  assign \$30  = \$33 ;
  assign \$35  = \$38 ;
  assign \$53  = \$54 ;
  assign \$52  = \$56 ;
  assign \$88  = \$89 ;
  assign rom_r_en = 1'h1;
  assign type_number = value[15:8];
  assign index = value[7:0];
  assign \$33  = { 2'h0, \$31 [32:2] };
  assign \$36  = { 2'h0, position_in_stream[5:2] };
endmodule
module handshake_detector(rx_valid, ack, nak, stall, nyet, usb_rst, usb_clk, rx_active, rx_data);
  reg \$auto$verilog_backend.cc:2083:dump_module$16  = 0;
  wire \$1 ;
  wire \$11 ;
  wire \$13 ;
  wire \$15 ;
  wire \$17 ;
  wire [3:0] \$19 ;
  wire \$21 ;
  wire \$23 ;
  wire \$25 ;
  wire \$27 ;
  wire [3:0] \$29 ;
  wire \$3 ;
  wire \$31 ;
  wire \$5 ;
  wire \$7 ;
  wire \$9 ;
  output ack;
  reg ack = 1'h0;
  reg \ack$next ;
  reg [3:0] active_pid = 4'h0;
  reg [3:0] \active_pid$next ;
  reg [1:0] fsm_state = 2'h0;
  reg [1:0] \fsm_state$next ;
  output nak;
  reg nak = 1'h0;
  reg \nak$next ;
  output nyet;
  reg nyet = 1'h0;
  reg \nyet$next ;
  input rx_active;
  wire rx_active;
  input [7:0] rx_data;
  wire [7:0] rx_data;
  input rx_valid;
  wire rx_valid;
  output stall;
  reg stall = 1'h0;
  reg \stall$next ;
  input usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  assign \$9  = ~  rx_active;
  assign \$11  = active_pid ==  4'he;
  assign \$13  = ~  rx_active;
  assign \$15  = active_pid ==  3'h6;
  assign \$17  = ~  rx_active;
  assign \$1  = ~  rx_active;
  assign \$19  = ~  rx_data[7:4];
  assign \$21  = rx_data[3:0] ==  \$19 ;
  assign \$23  = ~  rx_active;
  assign \$25  = ~  rx_active;
  assign \$27  = ~  rx_active;
  assign \$29  = ~  rx_data[7:4];
  assign \$31  = rx_data[3:0] ==  \$29 ;
  always @(posedge usb_clk)
    ack <= \ack$next ;
  always @(posedge usb_clk)
    nak <= \nak$next ;
  always @(posedge usb_clk)
    stall <= \stall$next ;
  always @(posedge usb_clk)
    nyet <= \nyet$next ;
  always @(posedge usb_clk)
    fsm_state <= \fsm_state$next ;
  always @(posedge usb_clk)
    active_pid <= \active_pid$next ;
  assign \$3  = active_pid ==  2'h2;
  assign \$5  = ~  rx_active;
  assign \$7  = active_pid ==  4'ha;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$16 ) begin end
    \ack$next  = 1'h0;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          ;
      2'h2:
          casez ({ rx_valid, \$1  })
            2'b?1:
                \ack$next  = \$3 ;
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \ack$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$16 ) begin end
    \nak$next  = 1'h0;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          ;
      2'h2:
          casez ({ rx_valid, \$5  })
            2'b?1:
                \nak$next  = \$7 ;
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \nak$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$16 ) begin end
    \stall$next  = 1'h0;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          ;
      2'h2:
          casez ({ rx_valid, \$9  })
            2'b?1:
                \stall$next  = \$11 ;
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \stall$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$16 ) begin end
    \nyet$next  = 1'h0;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          ;
      2'h2:
          casez ({ rx_valid, \$13  })
            2'b?1:
                \nyet$next  = \$15 ;
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \nyet$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$16 ) begin end
    \fsm_state$next  = fsm_state;
    casez (fsm_state)
      2'h0:
          casez (rx_active)
            1'h1:
                \fsm_state$next  = 2'h1;
          endcase
      2'h1:
          casez ({ rx_valid, \$17  })
            2'b?1:
                \fsm_state$next  = 2'h0;
            2'b1?:
                casez (\$21 )
                  1'h1:
                      \fsm_state$next  = 2'h2;
                  default:
                      \fsm_state$next  = 2'h3;
                endcase
          endcase
      2'h2:
          casez ({ rx_valid, \$23  })
            2'b?1:
                \fsm_state$next  = 2'h0;
            2'b1?:
                \fsm_state$next  = 2'h3;
          endcase
      2'h3:
          casez (\$25 )
            1'h1:
                \fsm_state$next  = 2'h0;
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \fsm_state$next  = 2'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$16 ) begin end
    \active_pid$next  = active_pid;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          casez ({ rx_valid, \$27  })
            2'b?1:
                ;
            2'b1?:
                casez (\$31 )
                  1'h1:
                      \active_pid$next  = rx_data[3:0];
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \active_pid$next  = 4'h0;
    endcase
  end
endmodule
module handshake_generator(issue_nak, issue_stall, usb_rst, usb_clk, valid, data, ready, issue_ack);
  reg \$auto$verilog_backend.cc:2083:dump_module$17  = 0;
  output [7:0] data;
  reg [7:0] data = 8'h00;
  reg [7:0] \data$next ;
  reg fsm_state = 1'h0;
  reg \fsm_state$next ;
  input issue_ack;
  wire issue_ack;
  input issue_nak;
  wire issue_nak;
  input issue_stall;
  wire issue_stall;
  input ready;
  wire ready;
  input usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  output valid;
  reg valid;
  always @(posedge usb_clk)
    data <= \data$next ;
  always @(posedge usb_clk)
    fsm_state <= \fsm_state$next ;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$17 ) begin end
    casez (fsm_state)
      1'h0:
          valid = 1'h0;
      1'h1:
          valid = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$17 ) begin end
    \data$next  = data;
    casez (fsm_state)
      1'h0:
        begin
          casez (issue_ack)
            1'h1:
                \data$next  = 8'hd2;
          endcase
          casez (issue_nak)
            1'h1:
                \data$next  = 8'h5a;
          endcase
          casez (issue_stall)
            1'h1:
                \data$next  = 8'h1e;
          endcase
        end
    endcase
    casez (usb_rst)
      1'h1:
          \data$next  = 8'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$17 ) begin end
    \fsm_state$next  = fsm_state;
    casez (fsm_state)
      1'h0:
        begin
          casez (issue_ack)
            1'h1:
                \fsm_state$next  = 1'h1;
          endcase
          casez (issue_nak)
            1'h1:
                \fsm_state$next  = 1'h1;
          endcase
          casez (issue_stall)
            1'h1:
                \fsm_state$next  = 1'h1;
          endcase
        end
      1'h1:
          casez (ready)
            1'h1:
                \fsm_state$next  = 1'h0;
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \fsm_state$next  = 1'h0;
    endcase
  end
endmodule
module receiver(rx_valid, valid, next, payload, packet_complete, crc_mismatch, ready_for_response, active_pid, usb_rst, usb_clk, rx_active, start, crc, \start$1 , tx_allowed, rx_data);
  reg \$auto$verilog_backend.cc:2083:dump_module$18  = 0;
  wire \$10 ;
  wire [3:0] \$12 ;
  wire \$14 ;
  wire \$16 ;
  wire \$18 ;
  wire \$2 ;
  wire \$20 ;
  wire \$22 ;
  wire \$24 ;
  wire \$26 ;
  wire \$28 ;
  wire \$30 ;
  wire [3:0] \$32 ;
  wire \$34 ;
  wire \$36 ;
  wire \$38 ;
  wire \$4 ;
  wire \$40 ;
  wire \$42 ;
  wire \$44 ;
  wire \$46 ;
  wire \$48 ;
  wire \$50 ;
  wire \$52 ;
  wire \$6 ;
  wire \$8 ;
  output [3:0] active_pid;
  reg [3:0] active_pid = 4'h0;
  reg [3:0] \active_pid$next ;
  input [15:0] crc;
  wire [15:0] crc;
  output crc_mismatch;
  reg crc_mismatch = 1'h0;
  reg \crc_mismatch$next ;
  reg [15:0] data_pipeline = 16'h0000;
  reg [15:0] \data_pipeline$next ;
  reg [2:0] fsm_state = 3'h0;
  reg [2:0] \fsm_state$next ;
  reg [15:0] last_byte_crc = 16'h0000;
  reg [15:0] \last_byte_crc$next ;
  reg [15:0] last_word_crc = 16'h0000;
  reg [15:0] \last_word_crc$next ;
  output next;
  reg next;
  output packet_complete;
  reg packet_complete = 1'h0;
  reg \packet_complete$next ;
  reg [3:0] packet_id = 4'h0;
  reg [3:0] \packet_id$next ;
  output [7:0] payload;
  reg [7:0] payload;
  output ready_for_response;
  reg ready_for_response;
  input rx_active;
  wire rx_active;
  input [7:0] rx_data;
  wire [7:0] rx_data;
  input rx_valid;
  wire rx_valid;
  output start;
  reg start;
  output \start$1 ;
  reg \start$1 ;
  input tx_allowed;
  wire tx_allowed;
  input usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  output valid;
  reg valid;
  assign \$10  = ~  rx_active;
  assign \$12  = ~  rx_data[7:4];
  assign \$14  = rx_data[3:0] ==  \$12 ;
  assign \$16  = rx_data[1:0] ==  2'h3;
  assign \$18  = \$14  &  \$16 ;
  assign \$20  = ~  rx_active;
  assign \$22  = ~  rx_active;
  assign \$24  = ~  rx_active;
  assign \$26  = last_word_crc ==  data_pipeline;
  assign \$28  = ~  rx_active;
  assign \$2  = ~  rx_active;
  assign \$30  = ~  rx_active;
  assign \$32  = ~  rx_data[7:4];
  assign \$34  = rx_data[3:0] ==  \$32 ;
  assign \$36  = rx_data[1:0] ==  2'h3;
  assign \$38  = \$34  &  \$36 ;
  assign \$40  = ~  rx_active;
  assign \$42  = ~  rx_active;
  assign \$44  = ~  rx_active;
  assign \$46  = ~  rx_active;
  assign \$48  = last_word_crc ==  data_pipeline;
  assign \$4  = last_word_crc ==  data_pipeline;
  assign \$50  = ~  rx_active;
  assign \$52  = last_word_crc ==  data_pipeline;
  always @(posedge usb_clk)
    packet_complete <= \packet_complete$next ;
  always @(posedge usb_clk)
    crc_mismatch <= \crc_mismatch$next ;
  always @(posedge usb_clk)
    fsm_state <= \fsm_state$next ;
  always @(posedge usb_clk)
    active_pid <= \active_pid$next ;
  always @(posedge usb_clk)
    data_pipeline <= \data_pipeline$next ;
  always @(posedge usb_clk)
    last_byte_crc <= \last_byte_crc$next ;
  always @(posedge usb_clk)
    last_word_crc <= \last_word_crc$next ;
  always @(posedge usb_clk)
    packet_id <= \packet_id$next ;
  assign \$6  = ~  rx_active;
  assign \$8  = last_word_crc ==  data_pipeline;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$18 ) begin end
    \packet_complete$next  = 1'h0;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          ;
      3'h4:
          ;
      3'h5:
          casez (\$2 )
            1'h1:
                casez (\$4 )
                  1'h1:
                      \packet_complete$next  = 1'h1;
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \packet_complete$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$18 ) begin end
    \crc_mismatch$next  = 1'h0;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          ;
      3'h4:
          ;
      3'h5:
          casez (\$6 )
            1'h1:
                casez (\$8 )
                  1'h1:
                      ;
                  default:
                      \crc_mismatch$next  = 1'h1;
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \crc_mismatch$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$18 ) begin end
    payload = 8'h00;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          ;
      3'h4:
          ;
      3'h5:
          casez (rx_valid)
            1'h1:
                payload = data_pipeline[7:0];
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$18 ) begin end
    \packet_id$next  = packet_id;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          ;
      3'h4:
          ;
      3'h5:
          casez (\$46 )
            1'h1:
                casez (\$48 )
                  1'h1:
                      \packet_id$next  = active_pid;
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \packet_id$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$18 ) begin end
    \start$1  = 1'h0;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          ;
      3'h4:
          ;
      3'h5:
          casez (\$50 )
            1'h1:
                casez (\$52 )
                  1'h1:
                      \start$1  = 1'h1;
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$18 ) begin end
    ready_for_response = 1'h0;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          ;
      3'h4:
          ;
      3'h5:
          ;
      3'h6:
          casez (tx_allowed)
            1'h1:
                ready_for_response = 1'h1;
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$18 ) begin end
    next = 1'h0;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          ;
      3'h4:
          ;
      3'h5:
          casez (rx_valid)
            1'h1:
                next = 1'h1;
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$18 ) begin end
    start = 1'h0;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          start = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$18 ) begin end
    \fsm_state$next  = fsm_state;
    casez (fsm_state)
      3'h0:
          casez (rx_active)
            1'h1:
                \fsm_state$next  = 3'h1;
          endcase
      3'h1:
          casez ({ rx_valid, \$10  })
            2'b?1:
                \fsm_state$next  = 3'h0;
            2'b1?:
                casez (\$18 )
                  1'h1:
                      \fsm_state$next  = 3'h2;
                  default:
                      \fsm_state$next  = 3'h3;
                endcase
          endcase
      3'h2:
        begin
          casez (rx_valid)
            1'h1:
                \fsm_state$next  = 3'h4;
          endcase
          casez (\$20 )
            1'h1:
                \fsm_state$next  = 3'h0;
          endcase
        end
      3'h4:
          casez ({ \$22 , rx_valid })
            2'b?1:
                \fsm_state$next  = 3'h5;
            2'b1?:
                \fsm_state$next  = 3'h0;
          endcase
      3'h5:
          casez (\$24 )
            1'h1:
                casez (\$26 )
                  1'h1:
                      \fsm_state$next  = 3'h6;
                  default:
                      \fsm_state$next  = 3'h0;
                endcase
          endcase
      3'h6:
          casez (tx_allowed)
            1'h1:
                \fsm_state$next  = 3'h0;
          endcase
      3'h3:
          casez (\$28 )
            1'h1:
                \fsm_state$next  = 3'h0;
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \fsm_state$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$18 ) begin end
    \active_pid$next  = active_pid;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          casez ({ rx_valid, \$30  })
            2'b?1:
                ;
            2'b1?:
                casez (\$38 )
                  1'h1:
                      \active_pid$next  = rx_data[3:0];
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \active_pid$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$18 ) begin end
    \data_pipeline$next  = data_pipeline;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          casez (rx_valid)
            1'h1:
                \data_pipeline$next [15:8] = rx_data;
          endcase
      3'h4:
          casez ({ \$40 , rx_valid })
            2'b?1:
              begin
                \data_pipeline$next [15:8] = rx_data;
                \data_pipeline$next [7:0] = data_pipeline[15:8];
              end
          endcase
      3'h5:
          casez (rx_valid)
            1'h1:
              begin
                \data_pipeline$next [15:8] = rx_data;
                \data_pipeline$next [7:0] = data_pipeline[15:8];
              end
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \data_pipeline$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$18 ) begin end
    \last_byte_crc$next  = last_byte_crc;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          casez (rx_valid)
            1'h1:
                \last_byte_crc$next  = crc;
          endcase
      3'h4:
          casez ({ \$42 , rx_valid })
            2'b?1:
                \last_byte_crc$next  = crc;
          endcase
      3'h5:
          casez (rx_valid)
            1'h1:
                \last_byte_crc$next  = crc;
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \last_byte_crc$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$18 ) begin end
    \last_word_crc$next  = last_word_crc;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          ;
      3'h4:
          casez ({ \$44 , rx_valid })
            2'b?1:
                \last_word_crc$next  = last_byte_crc;
          endcase
      3'h5:
          casez (rx_valid)
            1'h1:
                \last_word_crc$next  = last_byte_crc;
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \last_word_crc$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$18 ) begin end
    valid = 1'h0;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          ;
      3'h4:
          ;
      3'h5:
          valid = 1'h1;
    endcase
  end
endmodule
module register_window(usb_clk, busy, ulpi_data_in, ulpi_dir, ulpi_next, ulpi_data_out, ulpi_stop, done, address, write_data, read_request, write_request, usb_rst);
  reg \$auto$verilog_backend.cc:2083:dump_module$19  = 0;
  wire \$1 ;
  wire [7:0] \$11 ;
  wire \$13 ;
  wire [7:0] \$15 ;
  wire \$17 ;
  wire \$19 ;
  wire \$3 ;
  wire \$5 ;
  wire \$6 ;
  wire \$9 ;
  input [5:0] address;
  wire [5:0] address;
  output busy;
  wire busy;
  reg [5:0] current_address = 6'h00;
  reg [5:0] \current_address$next ;
  reg [7:0] current_write = 8'h00;
  reg [7:0] \current_write$next ;
  output done;
  reg done = 1'h0;
  reg \done$next ;
  reg [3:0] fsm_state = 4'h0;
  reg [3:0] \fsm_state$next ;
  reg [7:0] read_data = 8'h00;
  reg [7:0] \read_data$next ;
  input read_request;
  wire read_request;
  input [7:0] ulpi_data_in;
  wire [7:0] ulpi_data_in;
  output [7:0] ulpi_data_out;
  reg [7:0] ulpi_data_out = 8'h00;
  reg [7:0] \ulpi_data_out$next ;
  input ulpi_dir;
  wire ulpi_dir;
  input ulpi_next;
  wire ulpi_next;
  reg ulpi_out_req = 1'h0;
  reg \ulpi_out_req$next ;
  output ulpi_stop;
  reg ulpi_stop = 1'h0;
  reg \ulpi_stop$next ;
  input usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  input [7:0] write_data;
  wire [7:0] write_data;
  input write_request;
  wire write_request;
  assign \$9  = ~  ulpi_dir;
  assign \$11  = 8'hc0 |  address;
  assign \$13  = ~  ulpi_dir;
  assign \$15  = 8'h80 |  address;
  assign \$17  = ~  ulpi_dir;
  assign \$1  = ~  ulpi_dir;
  assign \$19  = ~  ulpi_dir;
  always @(posedge usb_clk)
    ulpi_out_req <= \ulpi_out_req$next ;
  always @(posedge usb_clk)
    ulpi_stop <= \ulpi_stop$next ;
  always @(posedge usb_clk)
    done <= \done$next ;
  always @(posedge usb_clk)
    ulpi_data_out <= \ulpi_data_out$next ;
  always @(posedge usb_clk)
    current_address <= \current_address$next ;
  always @(posedge usb_clk)
    current_write <= \current_write$next ;
  always @(posedge usb_clk)
    fsm_state <= \fsm_state$next ;
  always @(posedge usb_clk)
    read_data <= \read_data$next ;
  assign \$3  = ~  ulpi_dir;
  assign \$6  = !  fsm_state;
  assign \$5  = ~  \$6 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$19 ) begin end
    \ulpi_out_req$next  = 1'h0;
    casez (fsm_state)
      4'h0:
          ;
      4'h1:
          casez (\$1 )
            1'h1:
                \ulpi_out_req$next  = 1'h1;
          endcase
      4'h3:
        begin
          \ulpi_out_req$next  = 1'h1;
          casez ({ ulpi_next, ulpi_dir })
            2'b?1:
                \ulpi_out_req$next  = 1'h0;
            2'b1?:
                \ulpi_out_req$next  = 1'h0;
          endcase
        end
      4'h4:
          ;
      4'h5:
          ;
      4'h2:
          casez (\$3 )
            1'h1:
                \ulpi_out_req$next  = 1'h1;
          endcase
      4'h6:
        begin
          \ulpi_out_req$next  = 1'h1;
          casez ({ ulpi_next, ulpi_dir })
            2'b?1:
                \ulpi_out_req$next  = 1'h0;
          endcase
        end
      4'h7:
        begin
          \ulpi_out_req$next  = 1'h1;
          casez ({ ulpi_next, ulpi_dir })
            2'b?1:
                \ulpi_out_req$next  = 1'h0;
          endcase
        end
    endcase
    casez (usb_rst)
      1'h1:
          \ulpi_out_req$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$19 ) begin end
    \ulpi_stop$next  = 1'h0;
    casez (fsm_state)
      4'h0:
          ;
      4'h1:
          ;
      4'h3:
          ;
      4'h4:
          ;
      4'h5:
          ;
      4'h2:
          ;
      4'h6:
          ;
      4'h7:
          casez ({ ulpi_next, ulpi_dir })
            2'b?1:
                ;
            2'b1?:
                \ulpi_stop$next  = 1'h1;
          endcase
      4'h8:
          \ulpi_stop$next  = 1'h0;
    endcase
    casez (usb_rst)
      1'h1:
          \ulpi_stop$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$19 ) begin end
    \done$next  = 1'h0;
    casez (fsm_state)
      4'h0:
          ;
      4'h1:
          ;
      4'h3:
          ;
      4'h4:
          ;
      4'h5:
          \done$next  = 1'h1;
      4'h2:
          ;
      4'h6:
          ;
      4'h7:
          ;
      4'h8:
          \done$next  = 1'h1;
    endcase
    casez (usb_rst)
      1'h1:
          \done$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$19 ) begin end
    \ulpi_data_out$next  = ulpi_data_out;
    casez (fsm_state)
      4'h0:
          \ulpi_data_out$next  = 8'h00;
      4'h1:
          casez (\$9 )
            1'h1:
                \ulpi_data_out$next  = \$11 ;
          endcase
      4'h3:
          casez ({ ulpi_next, ulpi_dir })
            2'b?1:
                ;
            2'b1?:
                \ulpi_data_out$next  = 8'h00;
          endcase
      4'h4:
          ;
      4'h5:
          ;
      4'h2:
          casez (\$13 )
            1'h1:
                \ulpi_data_out$next  = \$15 ;
          endcase
      4'h6:
          casez ({ ulpi_next, ulpi_dir })
            2'b?1:
                ;
            2'b1?:
                \ulpi_data_out$next  = write_data;
          endcase
      4'h7:
          casez ({ ulpi_next, ulpi_dir })
            2'b?1:
                ;
            2'b1?:
                \ulpi_data_out$next  = 8'h00;
          endcase
      4'h8:
          \ulpi_data_out$next  = 8'h00;
    endcase
    casez (usb_rst)
      1'h1:
          \ulpi_data_out$next  = 8'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$19 ) begin end
    \current_address$next  = current_address;
    casez (fsm_state)
      4'h0:
          \current_address$next  = address;
    endcase
    casez (usb_rst)
      1'h1:
          \current_address$next  = 6'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$19 ) begin end
    \current_write$next  = current_write;
    casez (fsm_state)
      4'h0:
          \current_write$next  = write_data;
    endcase
    casez (usb_rst)
      1'h1:
          \current_write$next  = 8'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$19 ) begin end
    \fsm_state$next  = fsm_state;
    casez (fsm_state)
      4'h0:
        begin
          casez (read_request)
            1'h1:
                \fsm_state$next  = 4'h1;
          endcase
          casez (write_request)
            1'h1:
                \fsm_state$next  = 4'h2;
          endcase
        end
      4'h1:
          casez (\$17 )
            1'h1:
                \fsm_state$next  = 4'h3;
          endcase
      4'h3:
          casez ({ ulpi_next, ulpi_dir })
            2'b?1:
                \fsm_state$next  = 4'h1;
            2'b1?:
                \fsm_state$next  = 4'h4;
          endcase
      4'h4:
          \fsm_state$next  = 4'h5;
      4'h5:
          \fsm_state$next  = 4'h0;
      4'h2:
          casez (\$19 )
            1'h1:
                \fsm_state$next  = 4'h6;
          endcase
      4'h6:
          casez ({ ulpi_next, ulpi_dir })
            2'b?1:
                \fsm_state$next  = 4'h2;
            2'b1?:
                \fsm_state$next  = 4'h7;
          endcase
      4'h7:
          casez ({ ulpi_next, ulpi_dir })
            2'b?1:
                \fsm_state$next  = 4'h2;
            2'b1?:
                \fsm_state$next  = 4'h8;
          endcase
      4'h8:
          \fsm_state$next  = 4'h0;
    endcase
    casez (usb_rst)
      1'h1:
          \fsm_state$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$19 ) begin end
    \read_data$next  = read_data;
    casez (fsm_state)
      4'h0:
          ;
      4'h1:
          ;
      4'h3:
          ;
      4'h4:
          ;
      4'h5:
          \read_data$next  = ulpi_data_in;
    endcase
    casez (usb_rst)
      1'h1:
          \read_data$next  = 8'h00;
    endcase
  end
  assign busy = \$5 ;
endmodule
module request_mux(\type , is_in_request, request, value, index, length, received, pid, address, endpoint, new_token, ready_for_response, frame, new_frame, is_in, is_out, is_setup, is_ping, valid, first, last
, payload, ready, ack, nak, stall, \ack$1 , \nak$2 , \stall$3 , nyet, address_changed, new_address, active_config, config_changed, new_config, tx_data_pid, data_requested, \valid$4 , next, \payload$5 , rx_ready_for_response, status_requested
, \type$6 , \request$7 , \value$8 , \length$9 , \received$10 , \data_requested$11 , \status_requested$12 , \ack$13 , \active_config$14 , \type$15 , \request$16 , \data_requested$17 , \status_requested$18 , \rx_ready_for_response$19 , \type$20 , \data_requested$21 , \status_requested$22 , \address_changed$23 , \new_address$24 , \config_changed$25 , \new_config$26 
, \valid$27 , \tx_data_pid$28 , \valid$29 , \ack$30 , \ack$31 , \stall$32 , \stall$33 , \stall$34 , \payload$35 , \first$36 , \last$37 , \last$38 , \ready$39 , recipient);
  reg \$auto$verilog_backend.cc:2083:dump_module$20  = 0;
  wire \$124 ;
  wire \$127 ;
  wire \$131 ;
  wire \$134 ;
  wire \$136 ;
  wire \$138 ;
  output ack;
  wire ack;
  input \ack$1 ;
  wire \ack$1 ;
  wire \ack$105 ;
  wire \ack$126 ;
  output \ack$13 ;
  wire \ack$13 ;
  input \ack$30 ;
  wire \ack$30 ;
  input \ack$31 ;
  wire \ack$31 ;
  wire \ack$79 ;
  input [7:0] active_config;
  wire [7:0] active_config;
  wire [7:0] \active_config$109 ;
  output [7:0] \active_config$14 ;
  wire [7:0] \active_config$14 ;
  wire [7:0] \active_config$83 ;
  input [6:0] address;
  wire [6:0] address;
  wire [6:0] \address$45 ;
  wire [6:0] \address$69 ;
  wire [6:0] \address$95 ;
  output address_changed;
  reg address_changed;
  wire \address_changed$114 ;
  wire \address_changed$115 ;
  input \address_changed$23 ;
  wire \address_changed$23 ;
  output config_changed;
  reg config_changed;
  wire \config_changed$118 ;
  wire \config_changed$119 ;
  input \config_changed$25 ;
  wire \config_changed$25 ;
  input data_requested;
  wire data_requested;
  output \data_requested$11 ;
  wire \data_requested$11 ;
  output \data_requested$17 ;
  wire \data_requested$17 ;
  output \data_requested$21 ;
  wire \data_requested$21 ;
  input [3:0] endpoint;
  wire [3:0] endpoint;
  wire [3:0] \endpoint$46 ;
  wire [3:0] \endpoint$70 ;
  wire [3:0] \endpoint$96 ;
  output first;
  wire first;
  input \first$36 ;
  wire \first$36 ;
  input [10:0] frame;
  wire [10:0] frame;
  wire [10:0] \frame$49 ;
  wire [10:0] \frame$73 ;
  wire [10:0] \frame$99 ;
  input [15:0] index;
  wire [15:0] index;
  wire [15:0] \index$43 ;
  wire [15:0] \index$65 ;
  wire [15:0] \index$91 ;
  input is_in;
  wire is_in;
  wire \is_in$101 ;
  wire \is_in$51 ;
  wire \is_in$75 ;
  input is_in_request;
  wire is_in_request;
  wire \is_in_request$42 ;
  wire \is_in_request$63 ;
  wire \is_in_request$88 ;
  input is_out;
  wire is_out;
  wire \is_out$102 ;
  wire \is_out$52 ;
  wire \is_out$76 ;
  input is_ping;
  wire is_ping;
  wire \is_ping$104 ;
  wire \is_ping$54 ;
  wire \is_ping$78 ;
  input is_setup;
  wire is_setup;
  wire \is_setup$103 ;
  wire \is_setup$53 ;
  wire \is_setup$77 ;
  output last;
  wire last;
  input \last$37 ;
  wire \last$37 ;
  input \last$38 ;
  wire \last$38 ;
  input [15:0] length;
  wire [15:0] length;
  wire [15:0] \length$66 ;
  output [15:0] \length$9 ;
  wire [15:0] \length$9 ;
  wire [15:0] \length$92 ;
  output nak;
  wire nak;
  wire \nak$106 ;
  wire \nak$129 ;
  wire \nak$130 ;
  wire \nak$133 ;
  input \nak$2 ;
  wire \nak$2 ;
  wire \nak$55 ;
  wire \nak$80 ;
  output [6:0] new_address;
  reg [6:0] new_address;
  wire [6:0] \new_address$116 ;
  wire [6:0] \new_address$117 ;
  input [6:0] \new_address$24 ;
  wire [6:0] \new_address$24 ;
  output [7:0] new_config;
  reg [7:0] new_config;
  wire [7:0] \new_config$120 ;
  wire [7:0] \new_config$121 ;
  input [7:0] \new_config$26 ;
  wire [7:0] \new_config$26 ;
  input new_frame;
  wire new_frame;
  wire \new_frame$100 ;
  wire \new_frame$50 ;
  wire \new_frame$74 ;
  input new_token;
  wire new_token;
  wire \new_token$47 ;
  wire \new_token$71 ;
  wire \new_token$97 ;
  input next;
  wire next;
  wire \next$111 ;
  wire \next$59 ;
  wire \next$85 ;
  input nyet;
  wire nyet;
  wire \nyet$108 ;
  wire \nyet$57 ;
  wire \nyet$82 ;
  output [7:0] payload;
  wire [7:0] payload;
  wire [7:0] \payload$112 ;
  input [7:0] \payload$35 ;
  wire [7:0] \payload$35 ;
  input [7:0] \payload$5 ;
  wire [7:0] \payload$5 ;
  wire [7:0] \payload$60 ;
  wire [7:0] \payload$86 ;
  input [3:0] pid;
  wire [3:0] pid;
  wire [3:0] \pid$44 ;
  wire [3:0] \pid$68 ;
  wire [3:0] \pid$94 ;
  input ready;
  wire ready;
  output \ready$39 ;
  wire \ready$39 ;
  input ready_for_response;
  wire ready_for_response;
  wire \ready_for_response$48 ;
  wire \ready_for_response$72 ;
  wire \ready_for_response$98 ;
  input received;
  wire received;
  output \received$10 ;
  wire \received$10 ;
  wire \received$67 ;
  wire \received$93 ;
  input [4:0] recipient;
  wire [4:0] recipient;
  wire [4:0] \recipient$41 ;
  wire [4:0] \recipient$62 ;
  wire [4:0] \recipient$87 ;
  input [7:0] request;
  wire [7:0] request;
  output [7:0] \request$16 ;
  wire [7:0] \request$16 ;
  output [7:0] \request$7 ;
  wire [7:0] \request$7 ;
  wire [7:0] \request$89 ;
  input rx_ready_for_response;
  wire rx_ready_for_response;
  wire \rx_ready_for_response$113 ;
  output \rx_ready_for_response$19 ;
  wire \rx_ready_for_response$19 ;
  wire \rx_ready_for_response$61 ;
  output stall;
  wire stall;
  wire \stall$107 ;
  input \stall$3 ;
  wire \stall$3 ;
  input \stall$32 ;
  wire \stall$32 ;
  input \stall$33 ;
  wire \stall$33 ;
  input \stall$34 ;
  wire \stall$34 ;
  wire \stall$56 ;
  wire \stall$81 ;
  input status_requested;
  wire status_requested;
  output \status_requested$12 ;
  wire \status_requested$12 ;
  output \status_requested$18 ;
  wire \status_requested$18 ;
  output \status_requested$22 ;
  wire \status_requested$22 ;
  output tx_data_pid;
  reg tx_data_pid;
  wire \tx_data_pid$122 ;
  wire \tx_data_pid$123 ;
  input \tx_data_pid$28 ;
  wire \tx_data_pid$28 ;
  wire tx_mux_first;
  wire tx_mux_last;
  wire [7:0] tx_mux_payload;
  wire tx_mux_ready;
  wire tx_mux_valid;
  wire \tx_mux_valid$40 ;
  input [1:0] \type ;
  wire [1:0] \type ;
  output [1:0] \type$15 ;
  wire [1:0] \type$15 ;
  output [1:0] \type$20 ;
  wire [1:0] \type$20 ;
  output [1:0] \type$6 ;
  wire [1:0] \type$6 ;
  output valid;
  wire valid;
  wire \valid$110 ;
  input \valid$27 ;
  wire \valid$27 ;
  input \valid$29 ;
  wire \valid$29 ;
  input \valid$4 ;
  wire \valid$4 ;
  wire \valid$58 ;
  wire \valid$84 ;
  input [15:0] value;
  wire [15:0] value;
  wire [15:0] \value$64 ;
  output [15:0] \value$8 ;
  wire [15:0] \value$8 ;
  wire [15:0] \value$90 ;
  assign \$124  = \ack$30  |  \ack$31 ;
  assign \$136  = \stall$32  |  \stall$33 ;
  assign \$138  = \$136  |  \stall$34 ;
  \tx_mux$2  tx_mux (
    .first(tx_mux_first),
    .\first$5 (\first$36 ),
    .last(tx_mux_last),
    .\last$6 (\last$37 ),
    .\last$7 (\last$38 ),
    .payload(tx_mux_payload),
    .\payload$4 (\payload$35 ),
    .ready(tx_mux_ready),
    .\ready$8 (\ready$39 ),
    .valid(tx_mux_valid),
    .\valid$1 (\valid$27 ),
    .\valid$2 (\valid$29 ),
    .\valid$3 (1'h0)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$20 ) begin end
    address_changed = 1'h0;
    casez ({ \address_changed$115 , \address_changed$114 , \address_changed$23  })
      3'b??1:
          address_changed = \address_changed$23 ;
      3'b?1?:
          address_changed = 1'h0;
      3'b1??:
          address_changed = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$20 ) begin end
    new_address = 7'h00;
    casez ({ \address_changed$115 , \address_changed$114 , \address_changed$23  })
      3'b??1:
          new_address = \new_address$24 ;
      3'b?1?:
          new_address = 7'h00;
      3'b1??:
          new_address = 7'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$20 ) begin end
    config_changed = 1'h0;
    casez ({ \config_changed$119 , \config_changed$118 , \config_changed$25  })
      3'b??1:
          config_changed = \config_changed$25 ;
      3'b?1?:
          config_changed = 1'h0;
      3'b1??:
          config_changed = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$20 ) begin end
    new_config = 8'h00;
    casez ({ \config_changed$119 , \config_changed$118 , \config_changed$25  })
      3'b??1:
          new_config = \new_config$26 ;
      3'b?1?:
          new_config = 8'h00;
      3'b1??:
          new_config = 8'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$20 ) begin end
    tx_data_pid = 1'h1;
    casez (\valid$27 )
      1'h1:
          tx_data_pid = \tx_data_pid$28 ;
    endcase
    casez (\valid$29 )
      1'h1:
          tx_data_pid = 1'h1;
    endcase
    casez (\tx_mux_valid$40 )
      1'h1:
          tx_data_pid = 1'h1;
    endcase
  end
  assign \tx_mux_valid$40  = 1'h0;
  assign \address_changed$114  = 1'h0;
  assign \address_changed$115  = 1'h0;
  assign \new_address$116  = 7'h00;
  assign \new_address$117  = 7'h00;
  assign \config_changed$118  = 1'h0;
  assign \config_changed$119  = 1'h0;
  assign \new_config$120  = 8'h00;
  assign \new_config$121  = 8'h00;
  assign \tx_data_pid$122  = 1'h1;
  assign \tx_data_pid$123  = 1'h1;
  assign \ack$126  = 1'h0;
  assign \nak$129  = 1'h0;
  assign \nak$130  = 1'h0;
  assign \nak$133  = 1'h0;
  assign stall = \$138 ;
  assign nak = \$134 ;
  assign ack = \$127 ;
  assign tx_mux_ready = ready;
  assign payload = tx_mux_payload;
  assign last = tx_mux_last;
  assign first = tx_mux_first;
  assign valid = tx_mux_valid;
  assign \rx_ready_for_response$113  = rx_ready_for_response;
  assign \payload$112  = \payload$5 ;
  assign \next$111  = next;
  assign \valid$110  = \valid$4 ;
  assign \active_config$109  = active_config;
  assign \nyet$108  = nyet;
  assign \stall$107  = \stall$3 ;
  assign \nak$106  = \nak$2 ;
  assign \ack$105  = \ack$1 ;
  assign \status_requested$22  = status_requested;
  assign \data_requested$21  = data_requested;
  assign \is_ping$104  = is_ping;
  assign \is_setup$103  = is_setup;
  assign \is_out$102  = is_out;
  assign \is_in$101  = is_in;
  assign \new_frame$100  = new_frame;
  assign \frame$99  = frame;
  assign \ready_for_response$98  = ready_for_response;
  assign \new_token$97  = new_token;
  assign \endpoint$96  = endpoint;
  assign \address$95  = address;
  assign \pid$94  = pid;
  assign \received$93  = received;
  assign \length$92  = length;
  assign \index$91  = index;
  assign \value$90  = value;
  assign \request$89  = request;
  assign \is_in_request$88  = is_in_request;
  assign \type$20  = \type ;
  assign \recipient$87  = recipient;
  assign \rx_ready_for_response$19  = rx_ready_for_response;
  assign \payload$86  = \payload$5 ;
  assign \next$85  = next;
  assign \valid$84  = \valid$4 ;
  assign \active_config$83  = active_config;
  assign \nyet$82  = nyet;
  assign \stall$81  = \stall$3 ;
  assign \nak$80  = \nak$2 ;
  assign \ack$79  = \ack$1 ;
  assign \status_requested$18  = status_requested;
  assign \data_requested$17  = data_requested;
  assign \is_ping$78  = is_ping;
  assign \is_setup$77  = is_setup;
  assign \is_out$76  = is_out;
  assign \is_in$75  = is_in;
  assign \new_frame$74  = new_frame;
  assign \frame$73  = frame;
  assign \ready_for_response$72  = ready_for_response;
  assign \new_token$71  = new_token;
  assign \endpoint$70  = endpoint;
  assign \address$69  = address;
  assign \pid$68  = pid;
  assign \received$67  = received;
  assign \length$66  = length;
  assign \index$65  = index;
  assign \value$64  = value;
  assign \request$16  = request;
  assign \is_in_request$63  = is_in_request;
  assign \type$15  = \type ;
  assign \recipient$62  = recipient;
  assign \rx_ready_for_response$61  = rx_ready_for_response;
  assign \payload$60  = \payload$5 ;
  assign \next$59  = next;
  assign \valid$58  = \valid$4 ;
  assign \active_config$14  = active_config;
  assign \nyet$57  = nyet;
  assign \stall$56  = \stall$3 ;
  assign \nak$55  = \nak$2 ;
  assign \ack$13  = \ack$1 ;
  assign \status_requested$12  = status_requested;
  assign \data_requested$11  = data_requested;
  assign \is_ping$54  = is_ping;
  assign \is_setup$53  = is_setup;
  assign \is_out$52  = is_out;
  assign \is_in$51  = is_in;
  assign \new_frame$50  = new_frame;
  assign \frame$49  = frame;
  assign \ready_for_response$48  = ready_for_response;
  assign \new_token$47  = new_token;
  assign \endpoint$46  = endpoint;
  assign \address$45  = address;
  assign \pid$44  = pid;
  assign \received$10  = received;
  assign \length$9  = length;
  assign \index$43  = index;
  assign \value$8  = value;
  assign \request$7  = request;
  assign \is_in_request$42  = is_in_request;
  assign \type$6  = \type ;
  assign \recipient$41  = recipient;
  assign \$127  = \$124 ;
  assign \$131  = 1'h0;
  assign \$134  = 1'h0;
endmodule
module reset_sequencer(line_state, bus_reset, low_speed_only, full_speed_only, operating_mode, current_speed, termination_select, suspended, usb_rst, usb_clk, valid, data, bus_busy);
  reg \$auto$verilog_backend.cc:2083:dump_module$21  = 0;
  wire [18:0] \$1 ;
  wire \$10 ;
  wire \$101 ;
  wire \$103 ;
  wire \$105 ;
  wire \$107 ;
  wire \$109 ;
  wire \$111 ;
  wire \$113 ;
  wire \$115 ;
  wire \$117 ;
  wire \$119 ;
  wire \$12 ;
  wire \$121 ;
  wire \$123 ;
  wire \$125 ;
  wire \$127 ;
  wire \$129 ;
  wire \$131 ;
  wire \$133 ;
  wire \$135 ;
  wire \$137 ;
  wire \$139 ;
  wire \$14 ;
  wire \$141 ;
  wire \$143 ;
  wire \$145 ;
  wire \$147 ;
  wire \$149 ;
  wire \$151 ;
  wire \$153 ;
  wire \$155 ;
  wire \$157 ;
  wire \$159 ;
  wire \$16 ;
  wire \$161 ;
  wire \$163 ;
  wire \$165 ;
  wire \$167 ;
  wire [2:0] \$169 ;
  wire [2:0] \$170 ;
  wire \$18 ;
  wire [18:0] \$2 ;
  wire \$20 ;
  wire \$22 ;
  wire \$24 ;
  wire \$26 ;
  wire \$28 ;
  wire \$30 ;
  wire \$32 ;
  wire \$34 ;
  wire [18:0] \$36 ;
  wire [18:0] \$37 ;
  wire \$39 ;
  wire \$4 ;
  wire \$41 ;
  wire \$43 ;
  wire \$45 ;
  wire \$47 ;
  wire \$49 ;
  wire \$51 ;
  wire \$53 ;
  wire \$55 ;
  wire \$57 ;
  wire \$59 ;
  wire \$6 ;
  wire \$61 ;
  wire \$63 ;
  wire \$65 ;
  wire \$67 ;
  wire \$69 ;
  wire \$71 ;
  wire \$73 ;
  wire \$75 ;
  wire \$77 ;
  wire \$79 ;
  wire \$8 ;
  wire \$81 ;
  wire \$83 ;
  wire \$85 ;
  wire \$87 ;
  wire \$89 ;
  wire \$91 ;
  wire \$93 ;
  wire \$95 ;
  wire \$97 ;
  wire \$99 ;
  input bus_busy;
  wire bus_busy;
  reg bus_idle;
  output bus_reset;
  reg bus_reset;
  output [1:0] current_speed;
  reg [1:0] current_speed = 2'h1;
  reg [1:0] \current_speed$next ;
  output [7:0] data;
  reg [7:0] data;
  reg [3:0] fsm_state = 4'h0;
  reg [3:0] \fsm_state$next ;
  input full_speed_only;
  wire full_speed_only;
  input [1:0] line_state;
  wire [1:0] line_state;
  reg [17:0] line_state_time = 18'h00000;
  reg [17:0] \line_state_time$next ;
  input low_speed_only;
  wire low_speed_only;
  output [1:0] operating_mode;
  reg [1:0] operating_mode = 2'h0;
  reg [1:0] \operating_mode$next ;
  output suspended;
  reg suspended;
  output termination_select;
  reg termination_select = 1'h1;
  reg \termination_select$next ;
  reg [17:0] timer = 18'h00000;
  reg [17:0] \timer$next ;
  input usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  output valid;
  reg valid;
  reg [1:0] valid_pairs = 2'h0;
  reg [1:0] \valid_pairs$next ;
  reg was_hs_pre_suspend = 1'h0;
  reg \was_hs_pre_suspend$next ;
  assign \$99  = line_state ==  2'h2;
  assign \$101  = line_state_time ==  8'h96;
  assign \$103  = line_state !=  2'h2;
  assign \$105  = timer ==  18'h249f0;
  assign \$107  = timer ==  18'h249f0;
  assign \$10  = timer ==  18'h2bf20;
  assign \$109  = line_state ==  1'h1;
  assign \$111  = line_state_time ==  8'h96;
  assign \$113  = valid_pairs ==  2'h2;
  assign \$115  = line_state !=  1'h1;
  assign \$117  = timer ==  18'h249f0;
  assign \$119  = |  line_state;
  assign \$121  = timer ==  14'h2ee0;
  assign \$123  = line_state ==  1'h1;
  assign \$125  = line_state ==  1'h1;
  assign \$127  = low_speed_only &  \$125 ;
  assign \$12  = timer ==  17'h1d4c0;
  assign \$129  = ~  low_speed_only;
  assign \$131  = line_state ==  2'h2;
  assign \$133  = \$129  &  \$131 ;
  assign \$135  = \$127  |  \$133 ;
  assign \$137  = timer ==  8'h96;
  assign \$139  = low_speed_only |  full_speed_only;
  assign \$143  = timer ==  9'h12c;
  assign \$147  = timer ==  14'h2ee0;
  assign \$14  = |  line_state;
  assign \$149  = line_state ==  1'h1;
  assign \$151  = timer ==  8'h96;
  assign \$153  = line_state_time ==  18'h2bf20;
  assign \$155  = timer ==  14'h2ee0;
  assign \$157  = line_state ==  1'h1;
  assign \$159  = timer ==  18'h2bf20;
  assign \$161  = timer ==  18'h2bf20;
  assign \$163  = timer ==  17'h1d4c0;
  assign \$165  = line_state_time ==  8'h96;
  assign \$167  = valid_pairs ==  2'h2;
  assign \$16  = timer ==  14'h2ee0;
  assign \$170  = valid_pairs +  1'h1;
  always @(posedge usb_clk)
    timer <= \timer$next ;
  always @(posedge usb_clk)
    line_state_time <= \line_state_time$next ;
  always @(posedge usb_clk)
    current_speed <= \current_speed$next ;
  always @(posedge usb_clk)
    fsm_state <= \fsm_state$next ;
  always @(posedge usb_clk)
    was_hs_pre_suspend <= \was_hs_pre_suspend$next ;
  always @(posedge usb_clk)
    operating_mode <= \operating_mode$next ;
  always @(posedge usb_clk)
    termination_select <= \termination_select$next ;
  always @(posedge usb_clk)
    valid_pairs <= \valid_pairs$next ;
  assign \$18  = line_state ==  1'h1;
  assign \$20  = low_speed_only &  \$18 ;
  assign \$22  = ~  low_speed_only;
  assign \$24  = line_state ==  2'h2;
  assign \$26  = \$22  &  \$24 ;
  assign \$28  = \$20  |  \$26 ;
  assign \$2  = timer +  1'h1;
  assign \$30  = |  line_state;
  assign \$32  = timer ==  8'h96;
  assign \$34  = low_speed_only |  full_speed_only;
  assign \$37  = line_state_time +  1'h1;
  assign \$39  = ~  bus_idle;
  assign \$41  = line_state ==  2'h2;
  assign \$43  = line_state ==  1'h1;
  assign \$45  = |  line_state;
  assign \$47  = line_state ==  1'h1;
  assign \$4  = |  line_state;
  assign \$49  = low_speed_only &  \$47 ;
  assign \$51  = ~  low_speed_only;
  assign \$53  = line_state ==  2'h2;
  assign \$55  = \$51  &  \$53 ;
  assign \$57  = \$49  |  \$55 ;
  assign \$59  = timer ==  8'h96;
  assign \$61  = low_speed_only |  full_speed_only;
  assign \$63  = !  current_speed;
  assign \$65  = current_speed ==  1'h1;
  assign \$67  = !  line_state;
  assign \$69  = line_state ==  1'h1;
  assign \$71  = line_state ==  2'h2;
  assign \$73  = timer ==  18'h2bf20;
  assign \$75  = timer ==  9'h12c;
  assign \$77  = ~  low_speed_only;
  assign \$79  = ~  full_speed_only;
  assign \$81  = \$77  &  \$79 ;
  assign \$83  = line_state_time ==  18'h2bf20;
  assign \$87  = timer ==  18'h2bf20;
  assign \$8  = |  line_state;
  assign \$89  = full_speed_only |  low_speed_only;
  assign \$91  = ~  bus_busy;
  assign \$93  = ~  bus_busy;
  assign \$95  = timer ==  17'h1d4c0;
  assign \$97  = timer ==  18'h249f0;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$21 ) begin end
    \timer$next  = \$2 [17:0];
    casez (fsm_state)
      4'h0:
          \timer$next  = 18'h00000;
      4'h1:
        begin
          casez (\$4 )
            1'h1:
                \timer$next  = 18'h00000;
          endcase
          casez (\$6 )
            1'h1:
                \timer$next  = 18'h00000;
          endcase
        end
      4'h4:
        begin
          casez (\$8 )
            1'h1:
                \timer$next  = 18'h00000;
          endcase
          casez (\$10 )
            1'h1:
                \timer$next  = 18'h00000;
          endcase
        end
      4'h2:
          \timer$next  = 18'h00000;
      4'h7:
          ;
      4'h8:
          ;
      4'h9:
          casez (\$12 )
            1'h1:
                \timer$next  = 18'h00000;
          endcase
      4'ha:
          ;
      4'hb:
          ;
      4'hc:
          ;
      4'hd:
          ;
      4'he:
          \timer$next  = 18'h00000;
      4'h5:
          casez (\$14 )
            1'h1:
                \timer$next  = 18'h00000;
          endcase
      4'h6:
          casez (\$16 )
            1'h1:
                \timer$next  = 18'h00000;
          endcase
      4'h3:
        begin
          casez (\$28 )
            1'h1:
              begin
                \timer$next  = 18'h00000;
                casez (was_hs_pre_suspend)
                  1'h1:
                      ;
                  default:
                      \timer$next  = 18'h00000;
                endcase
              end
          endcase
          casez (\$30 )
            1'h1:
                \timer$next  = 18'h00000;
          endcase
          casez (\$32 )
            1'h1:
              begin
                \timer$next  = 18'h00000;
                casez (\$34 )
                  1'h1:
                      \timer$next  = 18'h00000;
                endcase
              end
          endcase
        end
    endcase
    casez (usb_rst)
      1'h1:
          \timer$next  = 18'h00000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$21 ) begin end
    \line_state_time$next  = \$37 [17:0];
    casez (fsm_state)
      4'h0:
          \line_state_time$next  = 18'h00000;
      4'h1:
          casez (\$39 )
            1'h1:
                \line_state_time$next  = 18'h00000;
          endcase
      4'h4:
          ;
      4'h2:
          ;
      4'h7:
          ;
      4'h8:
          ;
      4'h9:
          ;
      4'ha:
          casez (\$41 )
            1'h1:
                \line_state_time$next  = 18'h00000;
          endcase
      4'hb:
          ;
      4'hc:
          casez (\$43 )
            1'h1:
                \line_state_time$next  = 18'h00000;
          endcase
      4'hd:
          ;
      4'he:
          \line_state_time$next  = 18'h00000;
      4'h5:
          casez (\$45 )
            1'h1:
                \line_state_time$next  = 18'h00000;
          endcase
      4'h6:
          ;
      4'h3:
        begin
          casez (\$57 )
            1'h1:
                casez (was_hs_pre_suspend)
                  1'h1:
                      ;
                  default:
                      \line_state_time$next  = 18'h00000;
                endcase
          endcase
          casez (\$59 )
            1'h1:
                casez (\$61 )
                  1'h1:
                      \line_state_time$next  = 18'h00000;
                endcase
          endcase
        end
    endcase
    casez (usb_rst)
      1'h1:
          \line_state_time$next  = 18'h00000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$21 ) begin end
    data = 8'h00;
    casez (fsm_state)
      4'h0:
          ;
      4'h1:
          ;
      4'h4:
          ;
      4'h2:
          ;
      4'h7:
          ;
      4'h8:
          ;
      4'h9:
          data = 8'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$21 ) begin end
    \valid_pairs$next  = valid_pairs;
    casez (fsm_state)
      4'h0:
          ;
      4'h1:
          ;
      4'h4:
          ;
      4'h2:
          ;
      4'h7:
          ;
      4'h8:
          ;
      4'h9:
          casez (\$163 )
            1'h1:
                \valid_pairs$next  = 2'h0;
          endcase
      4'ha:
          ;
      4'hb:
          ;
      4'hc:
          ;
      4'hd:
          casez (\$165 )
            1'h1:
                casez (\$167 )
                  1'h1:
                      ;
                  default:
                      \valid_pairs$next  = \$170 [1:0];
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \valid_pairs$next  = 2'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$21 ) begin end
    suspended = 1'h0;
    casez (fsm_state)
      4'h0:
          ;
      4'h1:
          ;
      4'h4:
          ;
      4'h2:
          ;
      4'h7:
          ;
      4'h8:
          ;
      4'h9:
          ;
      4'ha:
          ;
      4'hb:
          ;
      4'hc:
          ;
      4'hd:
          ;
      4'he:
          ;
      4'h5:
          ;
      4'h6:
          ;
      4'h3:
          suspended = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$21 ) begin end
    casez ({ \$65 , \$63  })
      2'b?1:
          bus_idle = \$67 ;
      2'b1?:
          bus_idle = \$69 ;
      default:
          bus_idle = \$71 ;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$21 ) begin end
    \current_speed$next  = current_speed;
    casez (fsm_state)
      4'h0:
          casez (low_speed_only)
            1'h1:
                \current_speed$next  = 2'h2;
          endcase
      4'h1:
          ;
      4'h4:
          casez (\$73 )
            1'h1:
                \current_speed$next  = 2'h1;
          endcase
      4'h2:
          \current_speed$next  = 2'h0;
      4'h7:
          ;
      4'h8:
          ;
      4'h9:
          ;
      4'ha:
          ;
      4'hb:
          ;
      4'hc:
          ;
      4'hd:
          ;
      4'he:
          \current_speed$next  = 2'h0;
      4'h5:
          casez (low_speed_only)
            1'h1:
                \current_speed$next  = 2'h2;
            default:
                \current_speed$next  = 2'h1;
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \current_speed$next  = 2'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$21 ) begin end
    \fsm_state$next  = fsm_state;
    casez (fsm_state)
      4'h0:
          \fsm_state$next  = 4'h1;
      4'h1:
        begin
          casez (\$75 )
            1'h1:
                casez (\$81 )
                  1'h1:
                      \fsm_state$next  = 4'h2;
                endcase
          endcase
          casez (\$83 )
            1'h1:
                \fsm_state$next  = 4'h3;
          endcase
        end
      4'h4:
        begin
          casez (\$85 )
            1'h1:
                \fsm_state$next  = 4'h5;
          endcase
          casez (\$87 )
            1'h1:
                \fsm_state$next  = 4'h6;
          endcase
          casez (\$89 )
            1'h1:
                \fsm_state$next  = 4'h5;
          endcase
        end
      4'h2:
          \fsm_state$next  = 4'h7;
      4'h7:
          casez (\$91 )
            1'h1:
                \fsm_state$next  = 4'h8;
          endcase
      4'h8:
          casez (\$93 )
            1'h1:
                \fsm_state$next  = 4'h9;
          endcase
      4'h9:
          casez (\$95 )
            1'h1:
                \fsm_state$next  = 4'ha;
          endcase
      4'ha:
        begin
          casez (\$97 )
            1'h1:
                \fsm_state$next  = 4'h5;
          endcase
          casez (\$99 )
            1'h1:
                \fsm_state$next  = 4'hb;
          endcase
        end
      4'hb:
        begin
          casez (\$101 )
            1'h1:
                \fsm_state$next  = 4'hc;
          endcase
          casez (\$103 )
            1'h1:
                \fsm_state$next  = 4'ha;
          endcase
          casez (\$105 )
            1'h1:
                \fsm_state$next  = 4'h5;
          endcase
        end
      4'hc:
        begin
          casez (\$107 )
            1'h1:
                \fsm_state$next  = 4'h5;
          endcase
          casez (\$109 )
            1'h1:
                \fsm_state$next  = 4'hd;
          endcase
        end
      4'hd:
        begin
          casez (\$111 )
            1'h1:
                casez (\$113 )
                  1'h1:
                      \fsm_state$next  = 4'he;
                  default:
                      \fsm_state$next  = 4'ha;
                endcase
          endcase
          casez (\$115 )
            1'h1:
                \fsm_state$next  = 4'hc;
          endcase
          casez (\$117 )
            1'h1:
                \fsm_state$next  = 4'h5;
          endcase
        end
      4'he:
          \fsm_state$next  = 4'h4;
      4'h5:
          casez (\$119 )
            1'h1:
                \fsm_state$next  = 4'h1;
          endcase
      4'h6:
          casez (\$121 )
            1'h1:
                casez (\$123 )
                  1'h1:
                      \fsm_state$next  = 4'h3;
                  default:
                      \fsm_state$next  = 4'h2;
                endcase
          endcase
      4'h3:
        begin
          casez (\$135 )
            1'h1:
                casez (was_hs_pre_suspend)
                  1'h1:
                      \fsm_state$next  = 4'he;
                  default:
                      \fsm_state$next  = 4'h1;
                endcase
          endcase
          casez (\$137 )
            1'h1:
                casez (\$139 )
                  1'h1:
                      \fsm_state$next  = 4'h1;
                  default:
                      \fsm_state$next  = 4'h2;
                endcase
          endcase
        end
    endcase
    casez (usb_rst)
      1'h1:
          \fsm_state$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$21 ) begin end
    bus_reset = 1'h0;
    casez (fsm_state)
      4'h0:
          ;
      4'h1:
        begin
          casez (\$141 )
            1'h1:
                bus_reset = 1'h1;
          endcase
          casez (\$143 )
            1'h1:
                bus_reset = 1'h1;
          endcase
        end
      4'h4:
          casez (\$145 )
            1'h1:
                bus_reset = 1'h1;
          endcase
      4'h2:
          ;
      4'h7:
          ;
      4'h8:
          ;
      4'h9:
          ;
      4'ha:
          ;
      4'hb:
          ;
      4'hc:
          ;
      4'hd:
          ;
      4'he:
          ;
      4'h5:
          ;
      4'h6:
          casez (\$147 )
            1'h1:
                casez (\$149 )
                  1'h1:
                      ;
                  default:
                      bus_reset = 1'h1;
                endcase
          endcase
      4'h3:
          casez (\$151 )
            1'h1:
                bus_reset = 1'h1;
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$21 ) begin end
    \was_hs_pre_suspend$next  = was_hs_pre_suspend;
    casez (fsm_state)
      4'h0:
          ;
      4'h1:
          casez (\$153 )
            1'h1:
                \was_hs_pre_suspend$next  = 1'h0;
          endcase
      4'h4:
          ;
      4'h2:
          ;
      4'h7:
          ;
      4'h8:
          ;
      4'h9:
          ;
      4'ha:
          ;
      4'hb:
          ;
      4'hc:
          ;
      4'hd:
          ;
      4'he:
          ;
      4'h5:
          ;
      4'h6:
          casez (\$155 )
            1'h1:
                casez (\$157 )
                  1'h1:
                      \was_hs_pre_suspend$next  = 1'h1;
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \was_hs_pre_suspend$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$21 ) begin end
    \operating_mode$next  = operating_mode;
    casez (fsm_state)
      4'h0:
          ;
      4'h1:
          ;
      4'h4:
          casez (\$159 )
            1'h1:
                \operating_mode$next  = 2'h0;
          endcase
      4'h2:
          \operating_mode$next  = 2'h2;
      4'h7:
          ;
      4'h8:
          ;
      4'h9:
          ;
      4'ha:
          ;
      4'hb:
          ;
      4'hc:
          ;
      4'hd:
          ;
      4'he:
          \operating_mode$next  = 2'h0;
      4'h5:
          \operating_mode$next  = 2'h0;
    endcase
    casez (usb_rst)
      1'h1:
          \operating_mode$next  = 2'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$21 ) begin end
    \termination_select$next  = termination_select;
    casez (fsm_state)
      4'h0:
          ;
      4'h1:
          ;
      4'h4:
          casez (\$161 )
            1'h1:
                \termination_select$next  = 1'h1;
          endcase
      4'h2:
          \termination_select$next  = 1'h1;
      4'h7:
          ;
      4'h8:
          ;
      4'h9:
          ;
      4'ha:
          ;
      4'hb:
          ;
      4'hc:
          ;
      4'hd:
          ;
      4'he:
          \termination_select$next  = 1'h0;
      4'h5:
          \termination_select$next  = 1'h1;
    endcase
    casez (usb_rst)
      1'h1:
          \termination_select$next  = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$21 ) begin end
    valid = 1'h0;
    casez (fsm_state)
      4'h0:
          ;
      4'h1:
          ;
      4'h4:
          ;
      4'h2:
          ;
      4'h7:
          ;
      4'h8:
          ;
      4'h9:
          valid = 1'h1;
    endcase
  end
  assign \$1  = \$2 ;
  assign \$36  = \$37 ;
  assign \$169  = \$170 ;
  assign \$6  = 1'h0;
  assign \$85  = 1'h0;
  assign \$141  = 1'h0;
  assign \$145  = 1'h0;
endmodule
module rxevent_decoder(usb_clk, ulpi__dir__i, register_operation_in_progress, last_rx_command, ulpi__nxt, ulpi__data__i, line_state, vbus_valid, session_valid, session_end, rx_error, host_disconnect, id_digital, rx_stop, rx_start, usb_rst);
  reg \$auto$verilog_backend.cc:2083:dump_module$22  = 0;
  wire \$1 ;
  wire \$11 ;
  wire \$13 ;
  wire \$15 ;
  wire \$17 ;
  wire \$19 ;
  wire \$21 ;
  wire \$23 ;
  wire \$25 ;
  wire \$27 ;
  wire \$29 ;
  wire \$3 ;
  wire \$31 ;
  wire \$33 ;
  wire \$35 ;
  wire \$37 ;
  wire \$39 ;
  wire \$41 ;
  wire \$43 ;
  wire \$5 ;
  wire \$7 ;
  wire \$9 ;
  reg direction_delayed = 1'h0;
  reg \direction_delayed$next ;
  output host_disconnect;
  wire host_disconnect;
  output id_digital;
  wire id_digital;
  output [7:0] last_rx_command;
  reg [7:0] last_rx_command = 8'h00;
  reg [7:0] \last_rx_command$next ;
  output [1:0] line_state;
  wire [1:0] line_state;
  wire receiving;
  input register_operation_in_progress;
  wire register_operation_in_progress;
  wire rx_active;
  output rx_error;
  wire rx_error;
  output rx_start;
  reg rx_start = 1'h0;
  reg \rx_start$next ;
  output rx_stop;
  reg rx_stop = 1'h0;
  reg \rx_stop$next ;
  output session_end;
  wire session_end;
  output session_valid;
  wire session_valid;
  input [7:0] ulpi__data__i;
  wire [7:0] ulpi__data__i;
  input ulpi__dir__i;
  wire ulpi__dir__i;
  input ulpi__nxt;
  wire ulpi__nxt;
  input usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  output vbus_valid;
  wire vbus_valid;
  assign \$9  = \$5  &  \$7 ;
  assign \$11  = ~  rx_active;
  assign \$13  = \$11  &  ulpi__data__i[4];
  assign \$15  = ~  ulpi__nxt;
  assign \$17  = receiving &  \$15 ;
  assign \$1  = direction_delayed &  ulpi__dir__i;
  assign \$19  = ~  register_operation_in_progress;
  assign \$21  = \$17  &  \$19 ;
  assign \$23  = ~  ulpi__data__i[4];
  assign \$25  = rx_active &  \$23 ;
  assign \$27  = ~  ulpi__nxt;
  assign \$29  = receiving &  \$27 ;
  assign \$31  = ~  register_operation_in_progress;
  assign \$33  = \$29  &  \$31 ;
  assign \$35  = last_rx_command[3:2] ==  2'h3;
  assign \$37  = last_rx_command[3:2] ==  2'h2;
  assign \$3  = ~  ulpi__nxt;
  assign \$39  = !  last_rx_command[3:2];
  assign \$41  = last_rx_command[5:4] ==  2'h3;
  assign \$43  = last_rx_command[5:4] ==  2'h2;
  always @(posedge usb_clk)
    direction_delayed <= \direction_delayed$next ;
  always @(posedge usb_clk)
    rx_start <= \rx_start$next ;
  always @(posedge usb_clk)
    rx_stop <= \rx_stop$next ;
  always @(posedge usb_clk)
    last_rx_command <= \last_rx_command$next ;
  assign \$5  = receiving &  \$3 ;
  assign \$7  = ~  register_operation_in_progress;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$22 ) begin end
    \direction_delayed$next  = ulpi__dir__i;
    casez (usb_rst)
      1'h1:
          \direction_delayed$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$22 ) begin end
    \rx_start$next  = 1'h0;
    casez (\$9 )
      1'h1:
          casez (\$13 )
            1'h1:
                \rx_start$next  = 1'h1;
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \rx_start$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$22 ) begin end
    \rx_stop$next  = 1'h0;
    casez (\$21 )
      1'h1:
          casez (\$25 )
            1'h1:
                \rx_stop$next  = 1'h1;
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \rx_stop$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$22 ) begin end
    \last_rx_command$next  = last_rx_command;
    casez (\$33 )
      1'h1:
          \last_rx_command$next  = ulpi__data__i;
    endcase
    casez (usb_rst)
      1'h1:
          \last_rx_command$next  = 8'h00;
    endcase
  end
  assign id_digital = last_rx_command[6];
  assign host_disconnect = \$43 ;
  assign rx_error = \$41 ;
  assign rx_active = last_rx_command[4];
  assign session_end = \$39 ;
  assign session_valid = \$37 ;
  assign vbus_valid = \$35 ;
  assign line_state = last_rx_command[1:0];
  assign receiving = \$1 ;
endmodule
module setup_decoder(rx_valid, usb_rst, usb_clk, rx_active, start, crc, pid, new_token, speed, tx_allowed, \start$1 , recipient, \type , is_in_request, request, value, index, length, received, ack, rx_data
);
  reg \$auto$verilog_backend.cc:2083:dump_module$23  = 0;
  wire \$10 ;
  wire \$12 ;
  wire \$14 ;
  wire \$16 ;
  wire \$18 ;
  wire \$2 ;
  wire \$20 ;
  wire \$22 ;
  wire \$24 ;
  wire \$26 ;
  wire \$28 ;
  wire \$4 ;
  wire \$6 ;
  wire \$8 ;
  output ack;
  reg ack;
  input [15:0] crc;
  wire [15:0] crc;
  wire [15:0] data_handler_crc;
  wire [3:0] data_handler_length;
  wire data_handler_new_packet;
  wire [7:0] data_handler_packet_0;
  wire [7:0] data_handler_packet_1;
  wire [7:0] data_handler_packet_2;
  wire [7:0] data_handler_packet_3;
  wire [7:0] data_handler_packet_4;
  wire [7:0] data_handler_packet_5;
  wire [7:0] data_handler_packet_6;
  wire [7:0] data_handler_packet_7;
  wire data_handler_start;
  reg [1:0] fsm_state = 2'h0;
  reg [1:0] \fsm_state$next ;
  output [15:0] index;
  reg [15:0] index = 16'h0000;
  reg [15:0] \index$next ;
  output is_in_request;
  reg is_in_request = 1'h0;
  reg \is_in_request$next ;
  output [15:0] length;
  reg [15:0] length = 16'h0000;
  reg [15:0] \length$next ;
  input new_token;
  wire new_token;
  input [3:0] pid;
  wire [3:0] pid;
  output received;
  reg received = 1'h0;
  reg \received$next ;
  output [4:0] recipient;
  reg [4:0] recipient = 5'h00;
  reg [4:0] \recipient$next ;
  output [7:0] request;
  reg [7:0] request = 8'h00;
  reg [7:0] \request$next ;
  input rx_active;
  wire rx_active;
  input [7:0] rx_data;
  wire [7:0] rx_data;
  input rx_valid;
  wire rx_valid;
  input [1:0] speed;
  wire [1:0] speed;
  output start;
  wire start;
  output \start$1 ;
  wire \start$1 ;
  input tx_allowed;
  wire tx_allowed;
  output [1:0] \type ;
  reg [1:0] \type  = 2'h0;
  reg [1:0] \type$next ;
  input usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  output [15:0] value;
  reg [15:0] value = 16'h0000;
  reg [15:0] \value$next ;
  assign \$10  = !  speed;
  assign \$12  = tx_allowed |  \$10 ;
  assign \$14  = data_handler_length ==  4'h8;
  assign \$16  = data_handler_length ==  4'h8;
  assign \$18  = data_handler_length ==  4'h8;
  assign \$20  = data_handler_length ==  4'h8;
  assign \$22  = data_handler_length ==  4'h8;
  assign \$24  = data_handler_length ==  4'h8;
  assign \$26  = !  speed;
  assign \$28  = tx_allowed |  \$26 ;
  assign \$2  = data_handler_length ==  4'h8;
  always @(posedge usb_clk)
    received <= \received$next ;
  always @(posedge usb_clk)
    fsm_state <= \fsm_state$next ;
  always @(posedge usb_clk)
    recipient <= \recipient$next ;
  always @(posedge usb_clk)
    \type  <= \type$next ;
  always @(posedge usb_clk)
    is_in_request <= \is_in_request$next ;
  always @(posedge usb_clk)
    request <= \request$next ;
  always @(posedge usb_clk)
    value <= \value$next ;
  always @(posedge usb_clk)
    index <= \index$next ;
  always @(posedge usb_clk)
    length <= \length$next ;
  assign \$4  = pid ==  4'hd;
  assign \$6  = \$4  &  new_token;
  assign \$8  = data_handler_length ==  4'h8;
  data_handler data_handler (
    .crc(data_handler_crc),
    .length(data_handler_length),
    .new_packet(data_handler_new_packet),
    .packet_0(data_handler_packet_0),
    .packet_1(data_handler_packet_1),
    .packet_2(data_handler_packet_2),
    .packet_3(data_handler_packet_3),
    .packet_4(data_handler_packet_4),
    .packet_5(data_handler_packet_5),
    .packet_6(data_handler_packet_6),
    .packet_7(data_handler_packet_7),
    .rx_active(rx_active),
    .rx_data(rx_data),
    .rx_valid(rx_valid),
    .start(data_handler_start),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$23 ) begin end
    \index$next  = index;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          casez (data_handler_new_packet)
            1'h1:
                casez (\$20 )
                  1'h1:
                      \index$next  = { data_handler_packet_5, data_handler_packet_4 };
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \index$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$23 ) begin end
    \length$next  = length;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          casez (data_handler_new_packet)
            1'h1:
                casez (\$22 )
                  1'h1:
                      \length$next  = { data_handler_packet_7, data_handler_packet_6 };
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \length$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$23 ) begin end
    ack = 1'h0;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          casez (data_handler_new_packet)
            1'h1:
                casez (\$24 )
                  1'h1:
                      casez (\$28 )
                        1'h1:
                            ack = 1'h1;
                      endcase
                endcase
          endcase
      2'h2:
          casez (tx_allowed)
            1'h1:
                ack = 1'h1;
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$23 ) begin end
    \received$next  = 1'h0;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          casez (data_handler_new_packet)
            1'h1:
                casez (\$2 )
                  1'h1:
                      \received$next  = 1'h1;
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \received$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$23 ) begin end
    \fsm_state$next  = fsm_state;
    casez (fsm_state)
      2'h0:
          casez (\$6 )
            1'h1:
                \fsm_state$next  = 2'h1;
          endcase
      2'h1:
        begin
          casez (new_token)
            1'h1:
                \fsm_state$next  = 2'h0;
          endcase
          casez (data_handler_new_packet)
            1'h1:
                casez (\$8 )
                  1'h1:
                      casez (\$12 )
                        1'h1:
                            \fsm_state$next  = 2'h0;
                        default:
                            \fsm_state$next  = 2'h2;
                      endcase
                  default:
                      \fsm_state$next  = 2'h0;
                endcase
          endcase
        end
      2'h2:
          casez (tx_allowed)
            1'h1:
                \fsm_state$next  = 2'h0;
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \fsm_state$next  = 2'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$23 ) begin end
    \recipient$next  = recipient;
    \type$next  = \type ;
    \is_in_request$next  = is_in_request;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          casez (data_handler_new_packet)
            1'h1:
                casez (\$14 )
                  1'h1:
                      { \is_in_request$next , \type$next , \recipient$next  } = data_handler_packet_0;
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
        begin
          \recipient$next  = 5'h00;
          \type$next  = 2'h0;
          \is_in_request$next  = 1'h0;
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$23 ) begin end
    \request$next  = request;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          casez (data_handler_new_packet)
            1'h1:
                casez (\$16 )
                  1'h1:
                      \request$next  = data_handler_packet_1;
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \request$next  = 8'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$23 ) begin end
    \value$next  = value;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          casez (data_handler_new_packet)
            1'h1:
                casez (\$18 )
                  1'h1:
                      \value$next  = { data_handler_packet_3, data_handler_packet_2 };
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \value$next  = 16'h0000;
    endcase
  end
  assign \start$1  = data_handler_new_packet;
  assign data_handler_crc = crc;
  assign start = data_handler_start;
endmodule
module timer(usb_clk, speed, tx_allowed, start, usb_rst);
  reg \$auto$verilog_backend.cc:2083:dump_module$24  = 0;
  wire \$1 ;
  wire \$10 ;
  wire \$12 ;
  wire \$14 ;
  wire \$16 ;
  wire \$18 ;
  wire \$20 ;
  wire \$22 ;
  wire \$24 ;
  wire \$26 ;
  wire \$28 ;
  wire [10:0] \$3 ;
  wire \$30 ;
  wire \$32 ;
  wire \$34 ;
  wire [10:0] \$4 ;
  wire \$6 ;
  wire \$8 ;
  reg [9:0] counter = 10'h000;
  reg [9:0] \counter$next ;
  wire rx_timeout;
  reg rx_to_tx_at_max;
  reg rx_to_tx_at_min;
  input [1:0] speed;
  wire [1:0] speed;
  input start;
  wire start;
  output tx_allowed;
  wire tx_allowed;
  wire tx_timeout;
  reg tx_to_rx_timeout;
  input usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  assign \$10  = counter ==  1'h1;
  assign \$12  = counter ==  4'ha;
  assign \$14  = counter ==  1'h1;
  assign \$16  = !  speed;
  assign \$18  = speed ==  1'h1;
  assign \$1  = counter <  10'h281;
  assign \$20  = counter ==  5'h18;
  assign \$22  = counter ==  6'h20;
  assign \$24  = counter ==  5'h18;
  assign \$26  = !  speed;
  assign \$28  = speed ==  1'h1;
  assign \$30  = counter ==  7'h5c;
  assign \$32  = counter ==  7'h50;
  assign \$34  = counter ==  7'h5c;
  always @(posedge usb_clk)
    counter <= \counter$next ;
  assign \$4  = counter +  1'h1;
  assign \$6  = !  speed;
  assign \$8  = speed ==  1'h1;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$24 ) begin end
    \counter$next  = counter;
    casez ({ \$1 , start })
      2'b?1:
          \counter$next  = 10'h000;
      2'b1?:
          \counter$next  = \$4 [9:0];
    endcase
    casez (usb_rst)
      1'h1:
          \counter$next  = 10'h000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$24 ) begin end
    casez ({ \$8 , \$6  })
      2'b?1:
          rx_to_tx_at_min = \$10 ;
      2'b1?:
          rx_to_tx_at_min = \$12 ;
      default:
          rx_to_tx_at_min = \$14 ;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$24 ) begin end
    casez ({ \$18 , \$16  })
      2'b?1:
          rx_to_tx_at_max = \$20 ;
      2'b1?:
          rx_to_tx_at_max = \$22 ;
      default:
          rx_to_tx_at_max = \$24 ;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$24 ) begin end
    casez ({ \$28 , \$26  })
      2'b?1:
          tx_to_rx_timeout = \$30 ;
      2'b1?:
          tx_to_rx_timeout = \$32 ;
      default:
          tx_to_rx_timeout = \$34 ;
    endcase
  end
  assign \$3  = \$4 ;
  assign rx_timeout = tx_to_rx_timeout;
  assign tx_timeout = rx_to_tx_at_max;
  assign tx_allowed = rx_to_tx_at_min;
endmodule
module \timer$1 (usb_rst, usb_clk, start, tx_allowed, \start$1 , \tx_allowed$2 , tx_timeout, rx_timeout, speed);
  reg \$auto$verilog_backend.cc:2083:dump_module$25  = 0;
  wire \$10 ;
  wire \$12 ;
  wire \$14 ;
  wire \$16 ;
  wire \$18 ;
  wire \$20 ;
  wire \$22 ;
  wire \$24 ;
  wire \$26 ;
  wire \$28 ;
  wire \$3 ;
  wire \$30 ;
  wire \$32 ;
  wire \$34 ;
  wire \$36 ;
  wire \$38 ;
  wire \$5 ;
  wire [10:0] \$7 ;
  wire [10:0] \$8 ;
  reg [9:0] counter = 10'h000;
  reg [9:0] \counter$next ;
  output rx_timeout;
  wire rx_timeout;
  wire \rx_timeout$41 ;
  reg rx_to_tx_at_max;
  reg rx_to_tx_at_min;
  input [1:0] speed;
  wire [1:0] speed;
  input start;
  wire start;
  input \start$1 ;
  wire \start$1 ;
  output tx_allowed;
  wire tx_allowed;
  output \tx_allowed$2 ;
  wire \tx_allowed$2 ;
  output tx_timeout;
  wire tx_timeout;
  wire \tx_timeout$40 ;
  reg tx_to_rx_timeout;
  input usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  assign \$10  = !  speed;
  assign \$12  = speed ==  1'h1;
  assign \$14  = counter ==  1'h1;
  assign \$16  = counter ==  4'ha;
  assign \$18  = counter ==  1'h1;
  assign \$20  = !  speed;
  assign \$22  = speed ==  1'h1;
  assign \$24  = counter ==  5'h18;
  assign \$26  = counter ==  6'h20;
  assign \$28  = counter ==  5'h18;
  assign \$30  = !  speed;
  assign \$32  = speed ==  1'h1;
  assign \$34  = counter ==  7'h5c;
  assign \$36  = counter ==  7'h50;
  assign \$38  = counter ==  7'h5c;
  assign \$3  = start |  \start$1 ;
  always @(posedge usb_clk)
    counter <= \counter$next ;
  assign \$5  = counter <  10'h281;
  assign \$8  = counter +  1'h1;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$25 ) begin end
    \counter$next  = counter;
    casez ({ \$5 , \$3  })
      2'b?1:
          \counter$next  = 10'h000;
      2'b1?:
          \counter$next  = \$8 [9:0];
    endcase
    casez (usb_rst)
      1'h1:
          \counter$next  = 10'h000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$25 ) begin end
    casez ({ \$12 , \$10  })
      2'b?1:
          rx_to_tx_at_min = \$14 ;
      2'b1?:
          rx_to_tx_at_min = \$16 ;
      default:
          rx_to_tx_at_min = \$18 ;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$25 ) begin end
    casez ({ \$22 , \$20  })
      2'b?1:
          rx_to_tx_at_max = \$24 ;
      2'b1?:
          rx_to_tx_at_max = \$26 ;
      default:
          rx_to_tx_at_max = \$28 ;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$25 ) begin end
    casez ({ \$32 , \$30  })
      2'b?1:
          tx_to_rx_timeout = \$34 ;
      2'b1?:
          tx_to_rx_timeout = \$36 ;
      default:
          tx_to_rx_timeout = \$38 ;
    endcase
  end
  assign \$7  = \$8 ;
  assign rx_timeout = tx_to_rx_timeout;
  assign tx_timeout = rx_to_tx_at_max;
  assign \tx_allowed$2  = rx_to_tx_at_min;
  assign \rx_timeout$41  = tx_to_rx_timeout;
  assign \tx_timeout$40  = rx_to_tx_at_max;
  assign tx_allowed = rx_to_tx_at_min;
endmodule
module token_detector(rx_data, rx_valid, speed, pid, \address$1 , endpoint, new_token, ready_for_response, frame, new_frame, is_in, is_out, is_setup, is_ping, usb_rst, usb_clk, rx_active, address);
  reg \$auto$verilog_backend.cc:2083:dump_module$26  = 0;
  wire \$10 ;
  wire \$100 ;
  wire \$102 ;
  wire \$104 ;
  wire \$106 ;
  wire [3:0] \$108 ;
  wire \$110 ;
  wire \$112 ;
  wire \$114 ;
  wire [10:0] \$116 ;
  wire \$118 ;
  wire \$12 ;
  wire \$120 ;
  wire \$122 ;
  wire \$124 ;
  wire \$126 ;
  wire \$128 ;
  wire \$130 ;
  wire \$131 ;
  wire \$133 ;
  wire \$135 ;
  wire \$137 ;
  wire \$139 ;
  wire \$14 ;
  wire \$141 ;
  wire \$144 ;
  wire \$146 ;
  wire \$148 ;
  wire \$150 ;
  wire \$152 ;
  wire \$154 ;
  wire \$156 ;
  wire \$158 ;
  wire \$16 ;
  wire \$160 ;
  wire \$162 ;
  wire \$164 ;
  wire \$166 ;
  wire \$168 ;
  wire \$170 ;
  wire \$172 ;
  wire \$174 ;
  wire \$176 ;
  wire \$178 ;
  wire \$18 ;
  wire \$180 ;
  wire \$182 ;
  wire \$184 ;
  wire \$186 ;
  wire \$188 ;
  wire \$190 ;
  wire \$192 ;
  wire \$194 ;
  wire \$196 ;
  wire \$198 ;
  wire \$2 ;
  wire \$20 ;
  wire \$22 ;
  wire \$24 ;
  wire \$26 ;
  wire [3:0] \$28 ;
  wire \$30 ;
  wire \$32 ;
  wire \$34 ;
  wire \$36 ;
  wire \$38 ;
  wire \$4 ;
  wire \$40 ;
  wire \$42 ;
  wire \$44 ;
  wire \$46 ;
  wire \$48 ;
  wire \$49 ;
  wire \$51 ;
  wire \$53 ;
  wire \$55 ;
  wire \$57 ;
  wire \$59 ;
  wire \$6 ;
  wire \$62 ;
  wire \$64 ;
  wire \$66 ;
  wire \$68 ;
  wire \$70 ;
  wire \$72 ;
  wire \$74 ;
  wire \$76 ;
  wire \$78 ;
  wire \$8 ;
  wire \$80 ;
  wire \$82 ;
  wire \$84 ;
  wire \$86 ;
  wire \$88 ;
  wire \$90 ;
  wire \$92 ;
  wire \$94 ;
  wire \$96 ;
  wire \$98 ;
  input [6:0] address;
  wire [6:0] address;
  output [6:0] \address$1 ;
  reg [6:0] \address$1  = 7'h00;
  reg [6:0] \address$1$next ;
  reg [3:0] current_pid = 4'h0;
  reg [3:0] \current_pid$next ;
  output [3:0] endpoint;
  reg [3:0] endpoint = 4'h0;
  reg [3:0] \endpoint$next ;
  output [10:0] frame;
  reg [10:0] frame = 11'h000;
  reg [10:0] \frame$next ;
  reg [2:0] fsm_state = 3'h0;
  reg [2:0] \fsm_state$next ;
  output is_in;
  wire is_in;
  output is_out;
  wire is_out;
  output is_ping;
  wire is_ping;
  output is_setup;
  wire is_setup;
  output new_frame;
  reg new_frame = 1'h0;
  reg \new_frame$next ;
  output new_token;
  reg new_token = 1'h0;
  reg \new_token$next ;
  output [3:0] pid;
  reg [3:0] pid = 4'h0;
  reg [3:0] \pid$next ;
  output ready_for_response;
  wire ready_for_response;
  input rx_active;
  wire rx_active;
  input [7:0] rx_data;
  wire [7:0] rx_data;
  input rx_valid;
  wire rx_valid;
  input [1:0] speed;
  wire [1:0] speed;
  wire [1:0] timer_speed;
  reg timer_start;
  wire timer_tx_allowed;
  reg [10:0] token_data = 11'h000;
  reg [10:0] \token_data$next ;
  input usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  assign \$100  = ~  rx_active;
  assign \$102  = rx_data[1:0] ==  1'h1;
  assign \$104  = rx_data[3:0] ==  3'h4;
  assign \$106  = \$102  |  \$104 ;
  assign \$108  = ~  rx_data[7:4];
  assign \$10  = ~  rx_active;
  assign \$110  = rx_data[3:0] ==  \$108 ;
  assign \$112  = \$106  &  \$110 ;
  assign \$114  = ~  rx_active;
  assign \$116  = +  rx_data;
  assign \$118  = ~  rx_active;
  assign \$120  = token_data[0] ^  token_data[1];
  assign \$122  = \$120  ^  token_data[2];
  assign \$124  = \$122  ^  token_data[5];
  assign \$126  = \$124  ^  token_data[6];
  assign \$128  = \$126  ^  rx_data[0];
  assign \$12  = current_pid ==  3'h5;
  assign \$131  = token_data[0] ^  token_data[1];
  assign \$133  = \$131  ^  token_data[2];
  assign \$135  = \$133  ^  token_data[3];
  assign \$137  = \$135  ^  token_data[6];
  assign \$139  = \$137  ^  token_data[7];
  assign \$141  = \$139  ^  rx_data[1];
  assign \$130  = ~  \$141 ;
  assign \$144  = token_data[0] ^  token_data[1];
  assign \$146  = \$144  ^  token_data[2];
  assign \$148  = \$146  ^  token_data[3];
  assign \$14  = ~  rx_active;
  assign \$150  = \$148  ^  token_data[4];
  assign \$152  = \$150  ^  token_data[7];
  assign \$154  = \$152  ^  rx_data[0];
  assign \$156  = \$154  ^  rx_data[2];
  assign \$158  = token_data[0] ^  token_data[3];
  assign \$160  = \$158  ^  token_data[4];
  assign \$162  = \$160  ^  token_data[6];
  assign \$164  = \$162  ^  rx_data[1];
  assign \$166  = token_data[0] ^  token_data[1];
  assign \$168  = \$166  ^  token_data[4];
  assign \$16  = current_pid ==  3'h5;
  assign \$170  = \$168  ^  token_data[5];
  assign \$172  = \$170  ^  token_data[7];
  assign \$174  = \$172  ^  rx_data[2];
  assign \$176  = rx_data[7:3] ==  { \$174 , \$164 , \$156 , \$130 , \$128  };
  assign \$178  = ~  rx_active;
  assign \$180  = current_pid ==  3'h5;
  assign \$182  = ~  rx_active;
  assign \$184  = current_pid ==  3'h5;
  assign \$186  = token_data[6:0] ==  address;
  assign \$188  = ~  rx_active;
  assign \$18  = token_data[6:0] ==  address;
  assign \$190  = current_pid ==  3'h5;
  assign \$192  = token_data[6:0] ==  address;
  assign \$194  = ~  rx_active;
  assign \$196  = current_pid ==  3'h5;
  assign \$198  = token_data[6:0] ==  address;
  always @(posedge usb_clk)
    new_frame <= \new_frame$next ;
  always @(posedge usb_clk)
    new_token <= \new_token$next ;
  always @(posedge usb_clk)
    fsm_state <= \fsm_state$next ;
  always @(posedge usb_clk)
    current_pid <= \current_pid$next ;
  always @(posedge usb_clk)
    token_data <= \token_data$next ;
  always @(posedge usb_clk)
    frame <= \frame$next ;
  always @(posedge usb_clk)
    pid <= \pid$next ;
  always @(posedge usb_clk)
    \address$1  <= \address$1$next ;
  always @(posedge usb_clk)
    endpoint <= \endpoint$next ;
  assign \$20  = ~  rx_active;
  assign \$22  = rx_data[1:0] ==  1'h1;
  assign \$24  = rx_data[3:0] ==  3'h4;
  assign \$26  = \$22  |  \$24 ;
  assign \$28  = ~  rx_data[7:4];
  assign \$2  = pid ==  4'h9;
  assign \$30  = rx_data[3:0] ==  \$28 ;
  assign \$32  = \$26  &  \$30 ;
  assign \$34  = ~  rx_active;
  assign \$36  = ~  rx_active;
  assign \$38  = token_data[0] ^  token_data[1];
  assign \$40  = \$38  ^  token_data[2];
  assign \$42  = \$40  ^  token_data[5];
  assign \$44  = \$42  ^  token_data[6];
  assign \$46  = \$44  ^  rx_data[0];
  assign \$4  = pid ==  1'h1;
  assign \$49  = token_data[0] ^  token_data[1];
  assign \$51  = \$49  ^  token_data[2];
  assign \$53  = \$51  ^  token_data[3];
  assign \$55  = \$53  ^  token_data[6];
  assign \$57  = \$55  ^  token_data[7];
  assign \$59  = \$57  ^  rx_data[1];
  assign \$48  = ~  \$59 ;
  assign \$62  = token_data[0] ^  token_data[1];
  assign \$64  = \$62  ^  token_data[2];
  assign \$66  = \$64  ^  token_data[3];
  assign \$68  = \$66  ^  token_data[4];
  assign \$6  = pid ==  4'hd;
  assign \$70  = \$68  ^  token_data[7];
  assign \$72  = \$70  ^  rx_data[0];
  assign \$74  = \$72  ^  rx_data[2];
  assign \$76  = token_data[0] ^  token_data[3];
  assign \$78  = \$76  ^  token_data[4];
  assign \$80  = \$78  ^  token_data[6];
  assign \$82  = \$80  ^  rx_data[1];
  assign \$84  = token_data[0] ^  token_data[1];
  assign \$86  = \$84  ^  token_data[4];
  assign \$88  = \$86  ^  token_data[5];
  assign \$8  = pid ==  3'h4;
  assign \$90  = \$88  ^  token_data[7];
  assign \$92  = \$90  ^  rx_data[2];
  assign \$94  = rx_data[7:3] ==  { \$92 , \$82 , \$74 , \$48 , \$46  };
  assign \$96  = ~  rx_active;
  assign \$98  = ~  rx_active;
  timer timer (
    .speed(timer_speed),
    .start(timer_start),
    .tx_allowed(timer_tx_allowed),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$26 ) begin end
    \token_data$next  = token_data;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          casez ({ rx_valid, \$114  })
            2'b?1:
                ;
            2'b1?:
                \token_data$next  = \$116 ;
          endcase
      3'h4:
          casez ({ rx_valid, \$118  })
            2'b?1:
                ;
            2'b1?:
                casez (\$176 )
                  1'h1:
                      \token_data$next [10:8] = rx_data[2:0];
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \token_data$next  = 11'h000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$26 ) begin end
    \frame$next  = frame;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          ;
      3'h4:
          ;
      3'h5:
          casez ({ rx_valid, \$178  })
            2'b?1:
                casez (\$180 )
                  1'h1:
                      \frame$next  = token_data;
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \frame$next  = 11'h000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$26 ) begin end
    \pid$next  = pid;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          ;
      3'h4:
          ;
      3'h5:
          casez ({ rx_valid, \$182  })
            2'b?1:
                casez (\$184 )
                  1'h1:
                      ;
                  default:
                      casez (\$186 )
                        1'h1:
                            \pid$next  = current_pid;
                        default:
                            \pid$next  = 4'h0;
                      endcase
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \pid$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$26 ) begin end
    \address$1$next  = \address$1 ;
    \endpoint$next  = endpoint;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          ;
      3'h4:
          ;
      3'h5:
          casez ({ rx_valid, \$188  })
            2'b?1:
                casez (\$190 )
                  1'h1:
                      ;
                  default:
                      casez (\$192 )
                        1'h1:
                            { \endpoint$next , \address$1$next  } = token_data;
                      endcase
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
        begin
          \address$1$next  = 7'h00;
          \endpoint$next  = 4'h0;
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$26 ) begin end
    timer_start = 1'h0;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          ;
      3'h4:
          ;
      3'h5:
          casez ({ rx_valid, \$194  })
            2'b?1:
                casez (\$196 )
                  1'h1:
                      ;
                  default:
                      casez (\$198 )
                        1'h1:
                            timer_start = 1'h1;
                      endcase
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$26 ) begin end
    \new_frame$next  = 1'h0;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          ;
      3'h4:
          ;
      3'h5:
          casez ({ rx_valid, \$10  })
            2'b?1:
                casez (\$12 )
                  1'h1:
                      \new_frame$next  = 1'h1;
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \new_frame$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$26 ) begin end
    \new_token$next  = 1'h0;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h2:
          ;
      3'h4:
          ;
      3'h5:
          casez ({ rx_valid, \$14  })
            2'b?1:
                casez (\$16 )
                  1'h1:
                      ;
                  default:
                      casez (\$18 )
                        1'h1:
                            \new_token$next  = 1'h1;
                      endcase
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \new_token$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$26 ) begin end
    \fsm_state$next  = fsm_state;
    casez (fsm_state)
      3'h0:
          casez (rx_active)
            1'h1:
                \fsm_state$next  = 3'h1;
          endcase
      3'h1:
          casez ({ rx_valid, \$20  })
            2'b?1:
                \fsm_state$next  = 3'h0;
            2'b1?:
                casez (\$32 )
                  1'h1:
                      \fsm_state$next  = 3'h2;
                  default:
                      \fsm_state$next  = 3'h3;
                endcase
          endcase
      3'h2:
          casez ({ rx_valid, \$34  })
            2'b?1:
                \fsm_state$next  = 3'h0;
            2'b1?:
                \fsm_state$next  = 3'h4;
          endcase
      3'h4:
          casez ({ rx_valid, \$36  })
            2'b?1:
                \fsm_state$next  = 3'h0;
            2'b1?:
                casez (\$94 )
                  1'h1:
                      \fsm_state$next  = 3'h5;
                  default:
                      \fsm_state$next  = 3'h3;
                endcase
          endcase
      3'h5:
          casez ({ rx_valid, \$96  })
            2'b?1:
                \fsm_state$next  = 3'h0;
            2'b1?:
                \fsm_state$next  = 3'h3;
          endcase
      3'h3:
          casez (\$98 )
            1'h1:
                \fsm_state$next  = 3'h0;
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \fsm_state$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$26 ) begin end
    \current_pid$next  = current_pid;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          casez ({ rx_valid, \$100  })
            2'b?1:
                ;
            2'b1?:
                casez (\$112 )
                  1'h1:
                      \current_pid$next  = rx_data[3:0];
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \current_pid$next  = 4'h0;
    endcase
  end
  assign is_ping = \$8 ;
  assign is_setup = \$6 ;
  assign is_out = \$4 ;
  assign is_in = \$2 ;
  assign ready_for_response = timer_tx_allowed;
  assign timer_speed = speed;
endmodule
module translator(session_end, line_state, rx_data, rx_valid, tx_data, tx_valid, tx_ready, dm_pulldown, dp_pulldown, op_mode, xcvr_select, term_select, usb_rst, usb_clk, ulpi__clk, ulpi__rst, ulpi__data__oe, ulpi__dir__i, ulpi__nxt, ulpi__data__i, ulpi__data__o
, ulpi__stp, rx_active, busy);
  reg \$auto$verilog_backend.cc:2083:dump_module$27  = 0;
  wire \$1 ;
  wire \$11 ;
  wire \$13 ;
  wire \$15 ;
  wire \$17 ;
  wire \$19 ;
  wire \$21 ;
  wire \$23 ;
  wire \$25 ;
  wire \$27 ;
  wire \$29 ;
  wire \$3 ;
  wire \$5 ;
  wire \$7 ;
  wire \$9 ;
  reg \$sample$s$ulpi__dir__i$usb$1  = 1'h0;
  wire \$sample$s$ulpi__dir__i$usb$1$next ;
  output busy;
  wire busy;
  wire chrg_vbus;
  wire control_translator_bus_idle;
  wire control_translator_busy;
  wire control_translator_chrg_vbus;
  wire control_translator_dischrg_vbus;
  wire control_translator_dm_pulldown;
  wire control_translator_dp_pulldown;
  wire control_translator_id_pullup;
  wire [1:0] control_translator_op_mode;
  wire control_translator_suspend;
  wire control_translator_term_select;
  wire control_translator_use_external_vbus_indicator;
  wire [1:0] control_translator_xcvr_select;
  wire dischrg_vbus;
  input dm_pulldown;
  wire dm_pulldown;
  input dp_pulldown;
  wire dp_pulldown;
  wire host_disconnect;
  wire id_digital;
  wire id_pullup;
  wire [7:0] last_rx_command;
  output [1:0] line_state;
  wire [1:0] line_state;
  input [1:0] op_mode;
  wire [1:0] op_mode;
  wire [5:0] register_window_address;
  wire register_window_busy;
  wire register_window_done;
  wire register_window_read_request;
  wire [7:0] register_window_ulpi_data_in;
  wire [7:0] register_window_ulpi_data_out;
  wire register_window_ulpi_dir;
  wire register_window_ulpi_next;
  wire register_window_ulpi_stop;
  wire [7:0] register_window_write_data;
  wire register_window_write_request;
  output rx_active;
  reg rx_active = 1'h0;
  reg \rx_active$next ;
  output [7:0] rx_data;
  reg [7:0] rx_data = 8'h00;
  reg [7:0] \rx_data$next ;
  wire rx_error;
  output rx_valid;
  reg rx_valid = 1'h0;
  reg \rx_valid$next ;
  wire rxevent_decoder_host_disconnect;
  wire rxevent_decoder_id_digital;
  wire [7:0] rxevent_decoder_last_rx_command;
  wire [1:0] rxevent_decoder_line_state;
  wire rxevent_decoder_register_operation_in_progress;
  wire rxevent_decoder_rx_error;
  wire rxevent_decoder_rx_start;
  wire rxevent_decoder_rx_stop;
  wire rxevent_decoder_session_end;
  wire rxevent_decoder_session_valid;
  wire rxevent_decoder_vbus_valid;
  output session_end;
  wire session_end;
  wire session_valid;
  wire suspend;
  input term_select;
  wire term_select;
  wire transmit_translator_bus_idle;
  wire transmit_translator_busy;
  wire [1:0] transmit_translator_op_mode;
  wire [7:0] transmit_translator_tx_data;
  wire transmit_translator_tx_ready;
  wire transmit_translator_tx_valid;
  wire [7:0] transmit_translator_ulpi_data_out;
  wire transmit_translator_ulpi_nxt;
  wire transmit_translator_ulpi_out_req;
  wire transmit_translator_ulpi_stp;
  input [7:0] tx_data;
  wire [7:0] tx_data;
  output tx_ready;
  wire tx_ready;
  input tx_valid;
  wire tx_valid;
  input ulpi__clk;
  wire ulpi__clk;
  input [7:0] ulpi__data__i;
  wire [7:0] ulpi__data__i;
  output [7:0] ulpi__data__o;
  reg [7:0] ulpi__data__o;
  output ulpi__data__oe;
  wire ulpi__data__oe;
  input ulpi__dir__i;
  wire ulpi__dir__i;
  input ulpi__nxt;
  wire ulpi__nxt;
  output ulpi__rst;
  wire ulpi__rst;
  output ulpi__stp;
  reg ulpi__stp;
  output usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  wire use_external_vbus_indicator;
  wire vbus_valid;
  input [1:0] xcvr_select;
  wire [1:0] xcvr_select;
  assign \$9  = ~  control_translator_busy;
  assign \$11  = ~  ulpi__dir__i;
  assign \$13  = \$9  &  \$11 ;
  assign \$15  = ~  transmit_translator_busy;
  assign \$17  = ~  ulpi__dir__i;
  assign \$1  = ~  ulpi__dir__i;
  assign \$19  = \$17  |  rxevent_decoder_rx_stop;
  assign \$21  = ~  \$sample$s$ulpi__dir__i$usb$1 ;
  assign \$23  = \$21  &  ulpi__dir__i;
  assign \$25  = \$23  &  ulpi__nxt;
  assign \$27  = \$25  |  rxevent_decoder_rx_start;
  assign \$29  = ulpi__nxt &  rx_active;
  always @(posedge usb_clk)
    \$sample$s$ulpi__dir__i$usb$1  <= \$sample$s$ulpi__dir__i$usb$1$next ;
  always @(posedge usb_clk)
    rx_active <= \rx_active$next ;
  always @(posedge usb_clk)
    rx_data <= \rx_data$next ;
  always @(posedge usb_clk)
    rx_valid <= \rx_valid$next ;
  assign \$3  = register_window_busy |  transmit_translator_busy;
  assign \$5  = \$3  |  control_translator_busy;
  assign \$7  = \$5  |  ulpi__dir__i;
  control_translator control_translator (
    .address(register_window_address),
    .bus_idle(control_translator_bus_idle),
    .busy(register_window_busy),
    .\busy$1 (control_translator_busy),
    .chrg_vbus(1'h0),
    .dischrg_vbus(1'h0),
    .dm_pulldown(control_translator_dm_pulldown),
    .done(register_window_done),
    .dp_pulldown(control_translator_dp_pulldown),
    .id_pullup(1'h0),
    .op_mode(control_translator_op_mode),
    .read_request(register_window_read_request),
    .suspend(1'h0),
    .term_select(control_translator_term_select),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst),
    .use_external_vbus_indicator(1'h0),
    .write_data(register_window_write_data),
    .write_request(register_window_write_request),
    .xcvr_select(control_translator_xcvr_select)
  );
  register_window register_window (
    .address(register_window_address),
    .busy(register_window_busy),
    .done(register_window_done),
    .read_request(register_window_read_request),
    .ulpi_data_in(register_window_ulpi_data_in),
    .ulpi_data_out(register_window_ulpi_data_out),
    .ulpi_dir(register_window_ulpi_dir),
    .ulpi_next(register_window_ulpi_next),
    .ulpi_stop(register_window_ulpi_stop),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst),
    .write_data(register_window_write_data),
    .write_request(register_window_write_request)
  );
  rxevent_decoder rxevent_decoder (
    .host_disconnect(rxevent_decoder_host_disconnect),
    .id_digital(rxevent_decoder_id_digital),
    .last_rx_command(rxevent_decoder_last_rx_command),
    .line_state(rxevent_decoder_line_state),
    .register_operation_in_progress(rxevent_decoder_register_operation_in_progress),
    .rx_error(rxevent_decoder_rx_error),
    .rx_start(rxevent_decoder_rx_start),
    .rx_stop(rxevent_decoder_rx_stop),
    .session_end(rxevent_decoder_session_end),
    .session_valid(rxevent_decoder_session_valid),
    .ulpi__data__i(ulpi__data__i),
    .ulpi__dir__i(ulpi__dir__i),
    .ulpi__nxt(ulpi__nxt),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst),
    .vbus_valid(rxevent_decoder_vbus_valid)
  );
  transmit_translator transmit_translator (
    .bus_idle(transmit_translator_bus_idle),
    .busy(transmit_translator_busy),
    .op_mode(transmit_translator_op_mode),
    .tx_data(transmit_translator_tx_data),
    .tx_ready(transmit_translator_tx_ready),
    .tx_valid(transmit_translator_tx_valid),
    .ulpi_data_out(transmit_translator_ulpi_data_out),
    .ulpi_nxt(transmit_translator_ulpi_nxt),
    .ulpi_out_req(transmit_translator_ulpi_out_req),
    .ulpi_stp(transmit_translator_ulpi_stp),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$27 ) begin end
    casez (transmit_translator_ulpi_out_req)
      1'h1:
          ulpi__data__o = transmit_translator_ulpi_data_out;
      default:
          ulpi__data__o = register_window_ulpi_data_out;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$27 ) begin end
    casez (transmit_translator_ulpi_out_req)
      1'h1:
          ulpi__stp = transmit_translator_ulpi_stp;
      default:
          ulpi__stp = register_window_ulpi_stop;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$27 ) begin end
    \rx_active$next  = rx_active;
    casez ({ \$27 , \$19  })
      2'b?1:
          \rx_active$next  = 1'h0;
      2'b1?:
          \rx_active$next  = 1'h1;
    endcase
    casez (usb_rst)
      1'h1:
          \rx_active$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$27 ) begin end
    \rx_data$next  = ulpi__data__i;
    casez (usb_rst)
      1'h1:
          \rx_data$next  = 8'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$27 ) begin end
    \rx_valid$next  = \$29 ;
    casez (usb_rst)
      1'h1:
          \rx_valid$next  = 1'h0;
    endcase
  end
  assign suspend = 1'h0;
  assign id_pullup = 1'h0;
  assign chrg_vbus = 1'h0;
  assign dischrg_vbus = 1'h0;
  assign use_external_vbus_indicator = 1'h0;
  assign \$sample$s$ulpi__dir__i$usb$1$next  = ulpi__dir__i;
  assign control_translator_use_external_vbus_indicator = 1'h0;
  assign control_translator_dischrg_vbus = 1'h0;
  assign control_translator_chrg_vbus = 1'h0;
  assign control_translator_dp_pulldown = dp_pulldown;
  assign control_translator_dm_pulldown = dm_pulldown;
  assign control_translator_id_pullup = 1'h0;
  assign control_translator_suspend = 1'h0;
  assign control_translator_op_mode = op_mode;
  assign control_translator_term_select = term_select;
  assign control_translator_xcvr_select = xcvr_select;
  assign id_digital = rxevent_decoder_id_digital;
  assign host_disconnect = rxevent_decoder_host_disconnect;
  assign rx_error = rxevent_decoder_rx_error;
  assign session_end = rxevent_decoder_session_end;
  assign session_valid = rxevent_decoder_session_valid;
  assign vbus_valid = rxevent_decoder_vbus_valid;
  assign line_state = rxevent_decoder_line_state;
  assign register_window_ulpi_next = ulpi__nxt;
  assign register_window_ulpi_dir = ulpi__dir__i;
  assign register_window_ulpi_data_in = ulpi__data__i;
  assign control_translator_bus_idle = \$15 ;
  assign tx_ready = transmit_translator_tx_ready;
  assign transmit_translator_tx_valid = tx_valid;
  assign transmit_translator_tx_data = tx_data;
  assign transmit_translator_bus_idle = \$13 ;
  assign transmit_translator_op_mode = op_mode;
  assign transmit_translator_ulpi_nxt = ulpi__nxt;
  assign last_rx_command = rxevent_decoder_last_rx_command;
  assign rxevent_decoder_register_operation_in_progress = register_window_busy;
  assign busy = \$7 ;
  assign ulpi__data__oe = \$1 ;
  assign ulpi__rst = usb_rst;
  assign usb_clk = ulpi__clk;
endmodule
module transmit_translator(usb_clk, busy, ulpi_nxt, op_mode, bus_idle, tx_data, tx_valid, tx_ready, ulpi_out_req, ulpi_data_out, ulpi_stp, usb_rst);
  reg \$auto$verilog_backend.cc:2083:dump_module$28  = 0;
  wire \$1 ;
  wire \$11 ;
  wire \$13 ;
  wire \$15 ;
  wire [7:0] \$17 ;
  wire [6:0] \$18 ;
  wire \$2 ;
  wire \$21 ;
  wire \$23 ;
  wire \$25 ;
  wire \$27 ;
  wire \$29 ;
  wire \$5 ;
  wire \$7 ;
  wire \$9 ;
  input bus_idle;
  wire bus_idle;
  output busy;
  wire busy;
  reg fsm_state = 1'h0;
  reg \fsm_state$next ;
  input [1:0] op_mode;
  wire [1:0] op_mode;
  input [7:0] tx_data;
  wire [7:0] tx_data;
  output tx_ready;
  reg tx_ready;
  input tx_valid;
  wire tx_valid;
  output [7:0] ulpi_data_out;
  reg [7:0] ulpi_data_out;
  input ulpi_nxt;
  wire ulpi_nxt;
  output ulpi_out_req;
  reg ulpi_out_req = 1'h0;
  reg \ulpi_out_req$next ;
  output ulpi_stp;
  reg ulpi_stp;
  input usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  assign \$9  = op_mode ==  2'h2;
  assign \$11  = ~  tx_valid;
  assign \$13  = tx_valid &  bus_idle;
  assign \$15  = op_mode ==  2'h2;
  assign \$18  = 7'h40 |  tx_data[3:0];
  assign \$17  = +  \$18 ;
  assign \$21  = ~  tx_valid;
  assign \$23  = tx_valid &  bus_idle;
  assign \$25  = op_mode ==  2'h2;
  assign \$27  = tx_valid &  bus_idle;
  assign \$2  = ~  fsm_state;
  assign \$29  = ~  tx_valid;
  always @(posedge usb_clk)
    ulpi_out_req <= \ulpi_out_req$next ;
  always @(posedge usb_clk)
    fsm_state <= \fsm_state$next ;
  assign \$5  = ~  tx_valid;
  assign \$7  = tx_valid &  bus_idle;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$28 ) begin end
    casez (fsm_state)
      1'h0:
          ulpi_stp = 1'h0;
      1'h1:
        begin
          ulpi_stp = 1'h0;
          casez (\$5 )
            1'h1:
                ulpi_stp = 1'h1;
          endcase
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$28 ) begin end
    \ulpi_out_req$next  = ulpi_out_req;
    casez (fsm_state)
      1'h0:
          casez (\$7 )
            1'h1:
                casez (\$9 )
                  1'h1:
                      \ulpi_out_req$next  = 1'h1;
                  default:
                      \ulpi_out_req$next  = 1'h1;
                endcase
          endcase
      1'h1:
          casez (\$11 )
            1'h1:
                \ulpi_out_req$next  = 1'h0;
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \ulpi_out_req$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$28 ) begin end
    ulpi_data_out = 8'h00;
    casez (fsm_state)
      1'h0:
          casez (\$13 )
            1'h1:
                casez (\$15 )
                  1'h1:
                      ulpi_data_out = 8'h40;
                  default:
                      ulpi_data_out = \$17 ;
                endcase
          endcase
      1'h1:
        begin
          ulpi_data_out = tx_data;
          casez (\$21 )
            1'h1:
                ulpi_data_out = 8'h00;
          endcase
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$28 ) begin end
    tx_ready = 1'h0;
    casez (fsm_state)
      1'h0:
          casez (\$23 )
            1'h1:
                casez (\$25 )
                  1'h1:
                      tx_ready = 1'h0;
                  default:
                      tx_ready = ulpi_nxt;
                endcase
          endcase
      1'h1:
          tx_ready = ulpi_nxt;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$28 ) begin end
    \fsm_state$next  = fsm_state;
    casez (fsm_state)
      1'h0:
          casez (\$27 )
            1'h1:
                casez (ulpi_nxt)
                  1'h1:
                      \fsm_state$next  = 1'h1;
                endcase
          endcase
      1'h1:
          casez (\$29 )
            1'h1:
                \fsm_state$next  = 1'h0;
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \fsm_state$next  = 1'h0;
    endcase
  end
  assign busy = \$1 ;
  assign \$1  = fsm_state;
endmodule
module transmitter(first, last, payload, ready, data_pid, usb_rst, usb_clk, start, data, \valid$1 , \ready$2 , crc, valid);
  reg \$auto$verilog_backend.cc:2083:dump_module$29  = 0;
  wire \$11 ;
  wire \$13 ;
  wire \$15 ;
  wire \$3 ;
  wire \$5 ;
  wire \$7 ;
  wire \$9 ;
  input [15:0] crc;
  wire [15:0] crc;
  reg [7:0] current_data_pid = 8'h00;
  reg [7:0] \current_data_pid$next ;
  output [7:0] data;
  reg [7:0] data;
  input [1:0] data_pid;
  wire [1:0] data_pid;
  input first;
  wire first;
  reg [2:0] fsm_state = 3'h0;
  reg [2:0] \fsm_state$next ;
  reg is_zlp = 1'h0;
  reg \is_zlp$next ;
  input last;
  wire last;
  input [7:0] payload;
  wire [7:0] payload;
  output ready;
  reg ready;
  input \ready$2 ;
  wire \ready$2 ;
  reg [7:0] remaining_crc = 8'h00;
  reg [7:0] \remaining_crc$next ;
  output start;
  reg start;
  input usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  input valid;
  wire valid;
  output \valid$1 ;
  reg \valid$1 ;
  assign \$9  = last &  valid;
  assign \$11  = ~  valid;
  assign \$13  = last |  \$11 ;
  assign \$15  = \ready$2  &  \$13 ;
  always @(posedge usb_clk)
    current_data_pid <= \current_data_pid$next ;
  always @(posedge usb_clk)
    is_zlp <= \is_zlp$next ;
  always @(posedge usb_clk)
    fsm_state <= \fsm_state$next ;
  always @(posedge usb_clk)
    remaining_crc <= \remaining_crc$next ;
  assign \$3  = first &  valid;
  assign \$5  = last &  valid;
  assign \$7  = first &  valid;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$29 ) begin end
    ready = 1'h0;
    casez (fsm_state)
      3'h0:
          ready = 1'h0;
      3'h1:
          ready = 1'h0;
      3'h3:
          ready = \ready$2 ;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$29 ) begin end
    \current_data_pid$next  = current_data_pid;
    casez (fsm_state)
      3'h0:
          casez (data_pid)
            2'h0:
                \current_data_pid$next  = 8'hc3;
            2'h1:
                \current_data_pid$next  = 8'h4b;
            2'h2:
                \current_data_pid$next  = 8'h87;
            2'h?:
                \current_data_pid$next  = 8'h0f;
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \current_data_pid$next  = 8'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$29 ) begin end
    \is_zlp$next  = is_zlp;
    casez (fsm_state)
      3'h0:
          casez ({ \$5 , \$3  })
            2'b?1:
                \is_zlp$next  = 1'h0;
            2'b1?:
                \is_zlp$next  = 1'h1;
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \is_zlp$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$29 ) begin end
    \fsm_state$next  = fsm_state;
    casez (fsm_state)
      3'h0:
          casez ({ \$9 , \$7  })
            2'b?1:
                \fsm_state$next  = 3'h1;
            2'b1?:
                \fsm_state$next  = 3'h1;
          endcase
      3'h1:
          casez (\ready$2 )
            1'h1:
                casez (is_zlp)
                  1'h1:
                      \fsm_state$next  = 3'h2;
                  default:
                      \fsm_state$next  = 3'h3;
                endcase
          endcase
      3'h3:
          casez (\$15 )
            1'h1:
                \fsm_state$next  = 3'h2;
          endcase
      3'h2:
          casez (\ready$2 )
            1'h1:
                \fsm_state$next  = 3'h4;
          endcase
      3'h4:
          casez (\ready$2 )
            1'h1:
                \fsm_state$next  = 3'h0;
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \fsm_state$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$29 ) begin end
    start = 1'h0;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          start = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$29 ) begin end
    data = 8'h00;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          data = current_data_pid;
      3'h3:
          data = payload;
      3'h2:
          data = crc[7:0];
      3'h4:
          data = remaining_crc;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$29 ) begin end
    \valid$1  = 1'h0;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          \valid$1  = 1'h1;
      3'h3:
          \valid$1  = valid;
      3'h2:
          \valid$1  = 1'h1;
      3'h4:
          \valid$1  = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$29 ) begin end
    \remaining_crc$next  = remaining_crc;
    casez (fsm_state)
      3'h0:
          ;
      3'h1:
          ;
      3'h3:
          ;
      3'h2:
          \remaining_crc$next  = crc[15:8];
    endcase
    casez (usb_rst)
      1'h1:
          \remaining_crc$next  = 8'h00;
    endcase
  end
endmodule
module \transmitter$4 (usb_clk, valid, first, last, payload, ready, datum_0, datum_1, max_length, start, usb_rst);
  reg \$auto$verilog_backend.cc:2083:dump_module$30  = 0;
  wire \$1 ;
  wire \$11 ;
  wire \$13 ;
  wire \$15 ;
  wire [1:0] \$17 ;
  wire \$19 ;
  wire [1:0] \$21 ;
  wire \$23 ;
  wire \$25 ;
  wire [1:0] \$27 ;
  wire [1:0] \$28 ;
  wire \$3 ;
  wire \$30 ;
  wire \$32 ;
  wire [1:0] \$34 ;
  wire \$36 ;
  wire [1:0] \$38 ;
  wire \$40 ;
  wire \$42 ;
  wire \$5 ;
  wire [2:0] \$7 ;
  wire \$9 ;
  input [7:0] datum_0;
  wire [7:0] datum_0;
  input [7:0] datum_1;
  wire [7:0] datum_1;
  reg done;
  output first;
  wire first;
  reg [1:0] fsm_state = 2'h1;
  reg [1:0] \fsm_state$next ;
  output last;
  wire last;
  input [1:0] max_length;
  wire [1:0] max_length;
  output [7:0] payload;
  reg [7:0] payload;
  reg position_in_stream = 1'h0;
  reg \position_in_stream$next ;
  input ready;
  wire ready;
  input start;
  wire start;
  input usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  output valid;
  wire valid;
  assign \$9  = position_in_stream ==  \$7 ;
  assign \$11  = \$5  |  \$9 ;
  assign \$13  = \$11  &  valid;
  assign \$15  = !  fsm_state;
  assign \$17  = position_in_stream +  1'h1;
  assign \$1  = ~  position_in_stream;
  assign \$19  = \$17  <  max_length;
  assign \$21  = position_in_stream +  1'h1;
  assign \$23  = \$21  <  2'h2;
  assign \$25  = \$19  &  \$23 ;
  assign \$28  = position_in_stream +  1'h1;
  assign \$30  = max_length >  1'h0;
  assign \$32  = start &  \$30 ;
  assign \$34  = position_in_stream +  1'h1;
  assign \$36  = \$34  <  max_length;
  assign \$38  = position_in_stream +  1'h1;
  assign \$3  = \$1  &  valid;
  assign \$40  = \$38  <  2'h2;
  assign \$42  = \$36  &  \$40 ;
  always @(posedge usb_clk)
    position_in_stream <= \position_in_stream$next ;
  always @(posedge usb_clk)
    fsm_state <= \fsm_state$next ;
  assign \$7  = max_length -  1'h1;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$30 ) begin end
    \position_in_stream$next  = position_in_stream;
    casez (fsm_state)
      2'h1:
          \position_in_stream$next  = 1'h0;
      2'h0:
          casez (ready)
            1'h1:
                casez (\$25 )
                  1'h1:
                      \position_in_stream$next  = \$28 [0];
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \position_in_stream$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$30 ) begin end
    \fsm_state$next  = fsm_state;
    casez (fsm_state)
      2'h1:
          casez (\$32 )
            1'h1:
                \fsm_state$next  = 2'h0;
          endcase
      2'h0:
          casez (ready)
            1'h1:
                casez (\$42 )
                  1'h1:
                      ;
                  default:
                      \fsm_state$next  = 2'h2;
                endcase
          endcase
      2'h2:
          \fsm_state$next  = 2'h1;
    endcase
    casez (usb_rst)
      1'h1:
          \fsm_state$next  = 2'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$30 ) begin end
    payload = 8'h00;
    casez (fsm_state)
      2'h1:
          ;
      2'h0:
          casez (position_in_stream)
            1'h0:
                payload = datum_0;
            1'h?:
                payload = datum_1;
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$30 ) begin end
    done = 1'h0;
    casez (fsm_state)
      2'h1:
          ;
      2'h0:
          ;
      2'h2:
          done = 1'h1;
    endcase
  end
  assign \$27  = \$28 ;
  assign valid = \$15 ;
  assign last = \$13 ;
  assign first = \$3 ;
  assign \$5  = position_in_stream;
endmodule
module tx_manager(usb_clk, generate_zlps, active, valid, last, payload, ready, \valid$1 , first, \last$2 , \payload$3 , \ready$4 , data_pid, new_token, ready_for_response, is_in, nak, ack, usb_rst);
  reg \$auto$verilog_backend.cc:2083:dump_module$31  = 0;
  wire \$100 ;
  wire \$102 ;
  wire \$104 ;
  wire \$106 ;
  wire \$108 ;
  wire [10:0] \$11 ;
  wire \$110 ;
  wire \$112 ;
  wire [10:0] \$114 ;
  wire \$116 ;
  wire \$118 ;
  wire \$120 ;
  wire \$122 ;
  wire \$124 ;
  wire \$126 ;
  wire \$128 ;
  wire \$13 ;
  wire \$130 ;
  wire \$132 ;
  wire \$134 ;
  wire [10:0] \$136 ;
  wire \$138 ;
  wire \$140 ;
  wire \$142 ;
  wire \$144 ;
  wire \$146 ;
  wire \$148 ;
  wire \$15 ;
  wire [9:0] \$150 ;
  wire [9:0] \$151 ;
  wire [9:0] \$152 ;
  wire [9:0] \$153 ;
  wire [9:0] \$154 ;
  wire [9:0] \$155 ;
  wire \$156 ;
  wire [10:0] \$158 ;
  wire [10:0] \$159 ;
  wire \$161 ;
  wire [10:0] \$163 ;
  wire [10:0] \$164 ;
  wire [10:0] \$166 ;
  wire [10:0] \$167 ;
  wire \$169 ;
  wire \$17 ;
  wire \$171 ;
  wire \$173 ;
  wire \$175 ;
  wire \$177 ;
  wire \$179 ;
  wire \$181 ;
  wire \$183 ;
  wire \$185 ;
  wire \$187 ;
  wire [10:0] \$189 ;
  wire [10:0] \$19 ;
  wire [10:0] \$190 ;
  wire [10:0] \$192 ;
  wire [10:0] \$193 ;
  wire \$195 ;
  wire \$197 ;
  wire \$199 ;
  wire [10:0] \$201 ;
  wire \$203 ;
  wire \$205 ;
  wire \$207 ;
  wire [10:0] \$209 ;
  wire \$21 ;
  wire \$211 ;
  wire \$213 ;
  wire \$215 ;
  wire [10:0] \$217 ;
  wire \$219 ;
  wire \$221 ;
  wire \$223 ;
  wire [10:0] \$225 ;
  wire \$227 ;
  wire \$229 ;
  wire \$23 ;
  wire \$231 ;
  wire \$233 ;
  wire \$235 ;
  wire \$237 ;
  wire \$238 ;
  wire \$240 ;
  wire \$242 ;
  wire \$244 ;
  wire \$246 ;
  wire \$248 ;
  wire \$25 ;
  wire \$250 ;
  wire \$252 ;
  wire \$254 ;
  wire \$256 ;
  wire \$258 ;
  wire \$260 ;
  wire [10:0] \$262 ;
  wire \$264 ;
  wire \$266 ;
  wire \$268 ;
  wire \$270 ;
  wire \$272 ;
  wire \$274 ;
  wire \$276 ;
  wire \$278 ;
  wire [10:0] \$28 ;
  wire [10:0] \$280 ;
  wire \$282 ;
  wire \$284 ;
  wire \$286 ;
  wire \$288 ;
  wire \$290 ;
  wire \$292 ;
  wire \$294 ;
  wire \$296 ;
  wire \$298 ;
  wire \$30 ;
  wire \$300 ;
  wire \$302 ;
  wire \$304 ;
  wire [10:0] \$306 ;
  wire \$308 ;
  wire \$310 ;
  wire \$312 ;
  wire \$314 ;
  wire \$316 ;
  wire \$318 ;
  wire \$32 ;
  wire \$320 ;
  wire \$322 ;
  wire [10:0] \$324 ;
  wire \$326 ;
  wire \$328 ;
  wire \$330 ;
  wire \$332 ;
  wire \$334 ;
  wire \$336 ;
  wire [10:0] \$338 ;
  wire \$34 ;
  wire \$340 ;
  wire \$342 ;
  wire \$344 ;
  wire [10:0] \$346 ;
  wire \$348 ;
  wire \$350 ;
  wire [10:0] \$352 ;
  wire \$354 ;
  wire \$356 ;
  wire \$358 ;
  wire [10:0] \$36 ;
  wire [10:0] \$360 ;
  wire \$362 ;
  wire \$364 ;
  wire \$366 ;
  wire \$368 ;
  wire \$370 ;
  wire \$371 ;
  wire \$373 ;
  wire \$375 ;
  wire [10:0] \$377 ;
  wire \$379 ;
  wire \$38 ;
  wire [10:0] \$381 ;
  wire \$383 ;
  wire [10:0] \$385 ;
  wire \$387 ;
  wire \$389 ;
  wire \$391 ;
  wire \$393 ;
  wire \$395 ;
  wire \$397 ;
  wire \$399 ;
  wire \$40 ;
  wire \$401 ;
  wire \$403 ;
  wire \$405 ;
  wire [10:0] \$407 ;
  wire \$409 ;
  wire \$411 ;
  wire \$413 ;
  wire \$415 ;
  wire \$417 ;
  wire \$419 ;
  wire \$42 ;
  wire \$421 ;
  wire \$423 ;
  wire [10:0] \$425 ;
  wire \$427 ;
  wire \$429 ;
  wire \$431 ;
  wire \$433 ;
  wire \$435 ;
  wire \$437 ;
  wire \$439 ;
  wire \$44 ;
  wire \$441 ;
  wire \$443 ;
  wire \$445 ;
  wire \$447 ;
  wire \$449 ;
  wire [10:0] \$451 ;
  wire \$453 ;
  wire \$455 ;
  wire \$457 ;
  wire \$459 ;
  wire \$46 ;
  wire \$461 ;
  wire \$463 ;
  wire \$465 ;
  wire \$467 ;
  wire [10:0] \$469 ;
  wire \$471 ;
  wire \$473 ;
  wire \$475 ;
  wire \$477 ;
  wire [10:0] \$479 ;
  wire \$48 ;
  wire \$481 ;
  wire \$483 ;
  wire \$485 ;
  wire [10:0] \$487 ;
  wire \$489 ;
  wire \$491 ;
  wire \$493 ;
  wire [10:0] \$495 ;
  wire \$497 ;
  wire \$499 ;
  wire \$50 ;
  wire \$501 ;
  wire [10:0] \$503 ;
  wire \$505 ;
  wire \$507 ;
  wire \$509 ;
  wire \$511 ;
  wire \$513 ;
  wire \$515 ;
  wire \$517 ;
  wire \$519 ;
  wire \$52 ;
  wire \$521 ;
  wire \$523 ;
  wire \$525 ;
  wire \$527 ;
  wire [10:0] \$529 ;
  wire \$531 ;
  wire \$533 ;
  wire \$535 ;
  wire \$537 ;
  wire \$539 ;
  wire \$54 ;
  wire \$541 ;
  wire \$543 ;
  wire \$545 ;
  wire [10:0] \$547 ;
  wire \$549 ;
  wire \$551 ;
  wire \$553 ;
  wire \$555 ;
  wire \$557 ;
  wire \$559 ;
  wire \$56 ;
  wire \$561 ;
  wire \$563 ;
  wire \$565 ;
  wire \$567 ;
  wire \$569 ;
  wire \$571 ;
  wire [10:0] \$573 ;
  wire \$575 ;
  wire \$577 ;
  wire \$579 ;
  wire \$58 ;
  wire \$581 ;
  wire \$583 ;
  wire \$585 ;
  wire \$587 ;
  wire \$589 ;
  wire [10:0] \$591 ;
  wire \$593 ;
  wire \$595 ;
  wire \$597 ;
  wire \$599 ;
  wire \$60 ;
  wire [10:0] \$601 ;
  wire [10:0] \$602 ;
  wire \$604 ;
  wire \$606 ;
  wire \$608 ;
  wire \$609 ;
  wire \$611 ;
  wire \$613 ;
  wire \$615 ;
  wire \$617 ;
  wire \$619 ;
  wire [10:0] \$62 ;
  wire \$620 ;
  wire \$622 ;
  wire \$624 ;
  wire \$626 ;
  wire \$628 ;
  wire \$630 ;
  wire \$631 ;
  wire \$633 ;
  wire \$635 ;
  wire [10:0] \$637 ;
  wire \$639 ;
  wire \$64 ;
  wire [10:0] \$641 ;
  wire \$643 ;
  wire [10:0] \$645 ;
  wire \$647 ;
  wire \$66 ;
  wire \$68 ;
  wire [1:0] \$7 ;
  wire \$70 ;
  wire \$72 ;
  wire \$74 ;
  wire \$76 ;
  wire \$78 ;
  wire \$8 ;
  wire \$80 ;
  wire \$82 ;
  wire [10:0] \$84 ;
  wire \$86 ;
  wire \$88 ;
  wire \$90 ;
  wire \$92 ;
  wire \$94 ;
  wire \$96 ;
  wire \$98 ;
  reg [9:0] \$signal  = 10'h000;
  reg [9:0] \$signal$27  = 10'h000;
  reg [9:0] \$signal$27$next ;
  reg [9:0] \$signal$next ;
  input ack;
  wire ack;
  input active;
  wire active;
  reg buffer_toggle = 1'h0;
  reg \buffer_toggle$next ;
  output [1:0] data_pid;
  reg [1:0] data_pid = 2'h1;
  reg [1:0] \data_pid$next ;
  output first;
  reg first = 1'h0;
  reg \first$next ;
  reg [1:0] fsm_state = 2'h0;
  reg [1:0] \fsm_state$next ;
  input generate_zlps;
  wire generate_zlps;
  input is_in;
  wire is_in;
  input last;
  wire last;
  output \last$2 ;
  reg \last$2 ;
  output nak;
  reg nak;
  input new_token;
  wire new_token;
  input [7:0] payload;
  wire [7:0] payload;
  output [7:0] \payload$3 ;
  reg [7:0] \payload$3 ;
  output ready;
  reg ready;
  input \ready$4 ;
  wire \ready$4 ;
  input ready_for_response;
  wire ready_for_response;
  wire reset_sequence;
  reg [9:0] send_position = 10'h000;
  reg [9:0] \send_position$next ;
  wire start_with_data1;
  reg stream_ended_in_buffer0 = 1'h0;
  reg \stream_ended_in_buffer0$next ;
  reg stream_ended_in_buffer1 = 1'h0;
  reg \stream_ended_in_buffer1$next ;
  reg [8:0] transmit_buffer_0_r_addr;
  wire [7:0] transmit_buffer_0_r_data;
  reg [8:0] transmit_buffer_0_w_addr;
  wire [7:0] transmit_buffer_0_w_data;
  reg transmit_buffer_0_w_en;
  reg [8:0] transmit_buffer_1_r_addr;
  wire [7:0] transmit_buffer_1_r_data;
  reg [8:0] transmit_buffer_1_w_addr;
  wire [7:0] transmit_buffer_1_w_data;
  reg transmit_buffer_1_w_en;
  input usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  input valid;
  wire valid;
  output \valid$1 ;
  reg \valid$1 ;
  reg [7:0] transmit_buffer_0 [511:0];
  initial begin
    transmit_buffer_0[0] = 8'h00;
    transmit_buffer_0[1] = 8'h00;
    transmit_buffer_0[2] = 8'h00;
    transmit_buffer_0[3] = 8'h00;
    transmit_buffer_0[4] = 8'h00;
    transmit_buffer_0[5] = 8'h00;
    transmit_buffer_0[6] = 8'h00;
    transmit_buffer_0[7] = 8'h00;
    transmit_buffer_0[8] = 8'h00;
    transmit_buffer_0[9] = 8'h00;
    transmit_buffer_0[10] = 8'h00;
    transmit_buffer_0[11] = 8'h00;
    transmit_buffer_0[12] = 8'h00;
    transmit_buffer_0[13] = 8'h00;
    transmit_buffer_0[14] = 8'h00;
    transmit_buffer_0[15] = 8'h00;
    transmit_buffer_0[16] = 8'h00;
    transmit_buffer_0[17] = 8'h00;
    transmit_buffer_0[18] = 8'h00;
    transmit_buffer_0[19] = 8'h00;
    transmit_buffer_0[20] = 8'h00;
    transmit_buffer_0[21] = 8'h00;
    transmit_buffer_0[22] = 8'h00;
    transmit_buffer_0[23] = 8'h00;
    transmit_buffer_0[24] = 8'h00;
    transmit_buffer_0[25] = 8'h00;
    transmit_buffer_0[26] = 8'h00;
    transmit_buffer_0[27] = 8'h00;
    transmit_buffer_0[28] = 8'h00;
    transmit_buffer_0[29] = 8'h00;
    transmit_buffer_0[30] = 8'h00;
    transmit_buffer_0[31] = 8'h00;
    transmit_buffer_0[32] = 8'h00;
    transmit_buffer_0[33] = 8'h00;
    transmit_buffer_0[34] = 8'h00;
    transmit_buffer_0[35] = 8'h00;
    transmit_buffer_0[36] = 8'h00;
    transmit_buffer_0[37] = 8'h00;
    transmit_buffer_0[38] = 8'h00;
    transmit_buffer_0[39] = 8'h00;
    transmit_buffer_0[40] = 8'h00;
    transmit_buffer_0[41] = 8'h00;
    transmit_buffer_0[42] = 8'h00;
    transmit_buffer_0[43] = 8'h00;
    transmit_buffer_0[44] = 8'h00;
    transmit_buffer_0[45] = 8'h00;
    transmit_buffer_0[46] = 8'h00;
    transmit_buffer_0[47] = 8'h00;
    transmit_buffer_0[48] = 8'h00;
    transmit_buffer_0[49] = 8'h00;
    transmit_buffer_0[50] = 8'h00;
    transmit_buffer_0[51] = 8'h00;
    transmit_buffer_0[52] = 8'h00;
    transmit_buffer_0[53] = 8'h00;
    transmit_buffer_0[54] = 8'h00;
    transmit_buffer_0[55] = 8'h00;
    transmit_buffer_0[56] = 8'h00;
    transmit_buffer_0[57] = 8'h00;
    transmit_buffer_0[58] = 8'h00;
    transmit_buffer_0[59] = 8'h00;
    transmit_buffer_0[60] = 8'h00;
    transmit_buffer_0[61] = 8'h00;
    transmit_buffer_0[62] = 8'h00;
    transmit_buffer_0[63] = 8'h00;
    transmit_buffer_0[64] = 8'h00;
    transmit_buffer_0[65] = 8'h00;
    transmit_buffer_0[66] = 8'h00;
    transmit_buffer_0[67] = 8'h00;
    transmit_buffer_0[68] = 8'h00;
    transmit_buffer_0[69] = 8'h00;
    transmit_buffer_0[70] = 8'h00;
    transmit_buffer_0[71] = 8'h00;
    transmit_buffer_0[72] = 8'h00;
    transmit_buffer_0[73] = 8'h00;
    transmit_buffer_0[74] = 8'h00;
    transmit_buffer_0[75] = 8'h00;
    transmit_buffer_0[76] = 8'h00;
    transmit_buffer_0[77] = 8'h00;
    transmit_buffer_0[78] = 8'h00;
    transmit_buffer_0[79] = 8'h00;
    transmit_buffer_0[80] = 8'h00;
    transmit_buffer_0[81] = 8'h00;
    transmit_buffer_0[82] = 8'h00;
    transmit_buffer_0[83] = 8'h00;
    transmit_buffer_0[84] = 8'h00;
    transmit_buffer_0[85] = 8'h00;
    transmit_buffer_0[86] = 8'h00;
    transmit_buffer_0[87] = 8'h00;
    transmit_buffer_0[88] = 8'h00;
    transmit_buffer_0[89] = 8'h00;
    transmit_buffer_0[90] = 8'h00;
    transmit_buffer_0[91] = 8'h00;
    transmit_buffer_0[92] = 8'h00;
    transmit_buffer_0[93] = 8'h00;
    transmit_buffer_0[94] = 8'h00;
    transmit_buffer_0[95] = 8'h00;
    transmit_buffer_0[96] = 8'h00;
    transmit_buffer_0[97] = 8'h00;
    transmit_buffer_0[98] = 8'h00;
    transmit_buffer_0[99] = 8'h00;
    transmit_buffer_0[100] = 8'h00;
    transmit_buffer_0[101] = 8'h00;
    transmit_buffer_0[102] = 8'h00;
    transmit_buffer_0[103] = 8'h00;
    transmit_buffer_0[104] = 8'h00;
    transmit_buffer_0[105] = 8'h00;
    transmit_buffer_0[106] = 8'h00;
    transmit_buffer_0[107] = 8'h00;
    transmit_buffer_0[108] = 8'h00;
    transmit_buffer_0[109] = 8'h00;
    transmit_buffer_0[110] = 8'h00;
    transmit_buffer_0[111] = 8'h00;
    transmit_buffer_0[112] = 8'h00;
    transmit_buffer_0[113] = 8'h00;
    transmit_buffer_0[114] = 8'h00;
    transmit_buffer_0[115] = 8'h00;
    transmit_buffer_0[116] = 8'h00;
    transmit_buffer_0[117] = 8'h00;
    transmit_buffer_0[118] = 8'h00;
    transmit_buffer_0[119] = 8'h00;
    transmit_buffer_0[120] = 8'h00;
    transmit_buffer_0[121] = 8'h00;
    transmit_buffer_0[122] = 8'h00;
    transmit_buffer_0[123] = 8'h00;
    transmit_buffer_0[124] = 8'h00;
    transmit_buffer_0[125] = 8'h00;
    transmit_buffer_0[126] = 8'h00;
    transmit_buffer_0[127] = 8'h00;
    transmit_buffer_0[128] = 8'h00;
    transmit_buffer_0[129] = 8'h00;
    transmit_buffer_0[130] = 8'h00;
    transmit_buffer_0[131] = 8'h00;
    transmit_buffer_0[132] = 8'h00;
    transmit_buffer_0[133] = 8'h00;
    transmit_buffer_0[134] = 8'h00;
    transmit_buffer_0[135] = 8'h00;
    transmit_buffer_0[136] = 8'h00;
    transmit_buffer_0[137] = 8'h00;
    transmit_buffer_0[138] = 8'h00;
    transmit_buffer_0[139] = 8'h00;
    transmit_buffer_0[140] = 8'h00;
    transmit_buffer_0[141] = 8'h00;
    transmit_buffer_0[142] = 8'h00;
    transmit_buffer_0[143] = 8'h00;
    transmit_buffer_0[144] = 8'h00;
    transmit_buffer_0[145] = 8'h00;
    transmit_buffer_0[146] = 8'h00;
    transmit_buffer_0[147] = 8'h00;
    transmit_buffer_0[148] = 8'h00;
    transmit_buffer_0[149] = 8'h00;
    transmit_buffer_0[150] = 8'h00;
    transmit_buffer_0[151] = 8'h00;
    transmit_buffer_0[152] = 8'h00;
    transmit_buffer_0[153] = 8'h00;
    transmit_buffer_0[154] = 8'h00;
    transmit_buffer_0[155] = 8'h00;
    transmit_buffer_0[156] = 8'h00;
    transmit_buffer_0[157] = 8'h00;
    transmit_buffer_0[158] = 8'h00;
    transmit_buffer_0[159] = 8'h00;
    transmit_buffer_0[160] = 8'h00;
    transmit_buffer_0[161] = 8'h00;
    transmit_buffer_0[162] = 8'h00;
    transmit_buffer_0[163] = 8'h00;
    transmit_buffer_0[164] = 8'h00;
    transmit_buffer_0[165] = 8'h00;
    transmit_buffer_0[166] = 8'h00;
    transmit_buffer_0[167] = 8'h00;
    transmit_buffer_0[168] = 8'h00;
    transmit_buffer_0[169] = 8'h00;
    transmit_buffer_0[170] = 8'h00;
    transmit_buffer_0[171] = 8'h00;
    transmit_buffer_0[172] = 8'h00;
    transmit_buffer_0[173] = 8'h00;
    transmit_buffer_0[174] = 8'h00;
    transmit_buffer_0[175] = 8'h00;
    transmit_buffer_0[176] = 8'h00;
    transmit_buffer_0[177] = 8'h00;
    transmit_buffer_0[178] = 8'h00;
    transmit_buffer_0[179] = 8'h00;
    transmit_buffer_0[180] = 8'h00;
    transmit_buffer_0[181] = 8'h00;
    transmit_buffer_0[182] = 8'h00;
    transmit_buffer_0[183] = 8'h00;
    transmit_buffer_0[184] = 8'h00;
    transmit_buffer_0[185] = 8'h00;
    transmit_buffer_0[186] = 8'h00;
    transmit_buffer_0[187] = 8'h00;
    transmit_buffer_0[188] = 8'h00;
    transmit_buffer_0[189] = 8'h00;
    transmit_buffer_0[190] = 8'h00;
    transmit_buffer_0[191] = 8'h00;
    transmit_buffer_0[192] = 8'h00;
    transmit_buffer_0[193] = 8'h00;
    transmit_buffer_0[194] = 8'h00;
    transmit_buffer_0[195] = 8'h00;
    transmit_buffer_0[196] = 8'h00;
    transmit_buffer_0[197] = 8'h00;
    transmit_buffer_0[198] = 8'h00;
    transmit_buffer_0[199] = 8'h00;
    transmit_buffer_0[200] = 8'h00;
    transmit_buffer_0[201] = 8'h00;
    transmit_buffer_0[202] = 8'h00;
    transmit_buffer_0[203] = 8'h00;
    transmit_buffer_0[204] = 8'h00;
    transmit_buffer_0[205] = 8'h00;
    transmit_buffer_0[206] = 8'h00;
    transmit_buffer_0[207] = 8'h00;
    transmit_buffer_0[208] = 8'h00;
    transmit_buffer_0[209] = 8'h00;
    transmit_buffer_0[210] = 8'h00;
    transmit_buffer_0[211] = 8'h00;
    transmit_buffer_0[212] = 8'h00;
    transmit_buffer_0[213] = 8'h00;
    transmit_buffer_0[214] = 8'h00;
    transmit_buffer_0[215] = 8'h00;
    transmit_buffer_0[216] = 8'h00;
    transmit_buffer_0[217] = 8'h00;
    transmit_buffer_0[218] = 8'h00;
    transmit_buffer_0[219] = 8'h00;
    transmit_buffer_0[220] = 8'h00;
    transmit_buffer_0[221] = 8'h00;
    transmit_buffer_0[222] = 8'h00;
    transmit_buffer_0[223] = 8'h00;
    transmit_buffer_0[224] = 8'h00;
    transmit_buffer_0[225] = 8'h00;
    transmit_buffer_0[226] = 8'h00;
    transmit_buffer_0[227] = 8'h00;
    transmit_buffer_0[228] = 8'h00;
    transmit_buffer_0[229] = 8'h00;
    transmit_buffer_0[230] = 8'h00;
    transmit_buffer_0[231] = 8'h00;
    transmit_buffer_0[232] = 8'h00;
    transmit_buffer_0[233] = 8'h00;
    transmit_buffer_0[234] = 8'h00;
    transmit_buffer_0[235] = 8'h00;
    transmit_buffer_0[236] = 8'h00;
    transmit_buffer_0[237] = 8'h00;
    transmit_buffer_0[238] = 8'h00;
    transmit_buffer_0[239] = 8'h00;
    transmit_buffer_0[240] = 8'h00;
    transmit_buffer_0[241] = 8'h00;
    transmit_buffer_0[242] = 8'h00;
    transmit_buffer_0[243] = 8'h00;
    transmit_buffer_0[244] = 8'h00;
    transmit_buffer_0[245] = 8'h00;
    transmit_buffer_0[246] = 8'h00;
    transmit_buffer_0[247] = 8'h00;
    transmit_buffer_0[248] = 8'h00;
    transmit_buffer_0[249] = 8'h00;
    transmit_buffer_0[250] = 8'h00;
    transmit_buffer_0[251] = 8'h00;
    transmit_buffer_0[252] = 8'h00;
    transmit_buffer_0[253] = 8'h00;
    transmit_buffer_0[254] = 8'h00;
    transmit_buffer_0[255] = 8'h00;
    transmit_buffer_0[256] = 8'h00;
    transmit_buffer_0[257] = 8'h00;
    transmit_buffer_0[258] = 8'h00;
    transmit_buffer_0[259] = 8'h00;
    transmit_buffer_0[260] = 8'h00;
    transmit_buffer_0[261] = 8'h00;
    transmit_buffer_0[262] = 8'h00;
    transmit_buffer_0[263] = 8'h00;
    transmit_buffer_0[264] = 8'h00;
    transmit_buffer_0[265] = 8'h00;
    transmit_buffer_0[266] = 8'h00;
    transmit_buffer_0[267] = 8'h00;
    transmit_buffer_0[268] = 8'h00;
    transmit_buffer_0[269] = 8'h00;
    transmit_buffer_0[270] = 8'h00;
    transmit_buffer_0[271] = 8'h00;
    transmit_buffer_0[272] = 8'h00;
    transmit_buffer_0[273] = 8'h00;
    transmit_buffer_0[274] = 8'h00;
    transmit_buffer_0[275] = 8'h00;
    transmit_buffer_0[276] = 8'h00;
    transmit_buffer_0[277] = 8'h00;
    transmit_buffer_0[278] = 8'h00;
    transmit_buffer_0[279] = 8'h00;
    transmit_buffer_0[280] = 8'h00;
    transmit_buffer_0[281] = 8'h00;
    transmit_buffer_0[282] = 8'h00;
    transmit_buffer_0[283] = 8'h00;
    transmit_buffer_0[284] = 8'h00;
    transmit_buffer_0[285] = 8'h00;
    transmit_buffer_0[286] = 8'h00;
    transmit_buffer_0[287] = 8'h00;
    transmit_buffer_0[288] = 8'h00;
    transmit_buffer_0[289] = 8'h00;
    transmit_buffer_0[290] = 8'h00;
    transmit_buffer_0[291] = 8'h00;
    transmit_buffer_0[292] = 8'h00;
    transmit_buffer_0[293] = 8'h00;
    transmit_buffer_0[294] = 8'h00;
    transmit_buffer_0[295] = 8'h00;
    transmit_buffer_0[296] = 8'h00;
    transmit_buffer_0[297] = 8'h00;
    transmit_buffer_0[298] = 8'h00;
    transmit_buffer_0[299] = 8'h00;
    transmit_buffer_0[300] = 8'h00;
    transmit_buffer_0[301] = 8'h00;
    transmit_buffer_0[302] = 8'h00;
    transmit_buffer_0[303] = 8'h00;
    transmit_buffer_0[304] = 8'h00;
    transmit_buffer_0[305] = 8'h00;
    transmit_buffer_0[306] = 8'h00;
    transmit_buffer_0[307] = 8'h00;
    transmit_buffer_0[308] = 8'h00;
    transmit_buffer_0[309] = 8'h00;
    transmit_buffer_0[310] = 8'h00;
    transmit_buffer_0[311] = 8'h00;
    transmit_buffer_0[312] = 8'h00;
    transmit_buffer_0[313] = 8'h00;
    transmit_buffer_0[314] = 8'h00;
    transmit_buffer_0[315] = 8'h00;
    transmit_buffer_0[316] = 8'h00;
    transmit_buffer_0[317] = 8'h00;
    transmit_buffer_0[318] = 8'h00;
    transmit_buffer_0[319] = 8'h00;
    transmit_buffer_0[320] = 8'h00;
    transmit_buffer_0[321] = 8'h00;
    transmit_buffer_0[322] = 8'h00;
    transmit_buffer_0[323] = 8'h00;
    transmit_buffer_0[324] = 8'h00;
    transmit_buffer_0[325] = 8'h00;
    transmit_buffer_0[326] = 8'h00;
    transmit_buffer_0[327] = 8'h00;
    transmit_buffer_0[328] = 8'h00;
    transmit_buffer_0[329] = 8'h00;
    transmit_buffer_0[330] = 8'h00;
    transmit_buffer_0[331] = 8'h00;
    transmit_buffer_0[332] = 8'h00;
    transmit_buffer_0[333] = 8'h00;
    transmit_buffer_0[334] = 8'h00;
    transmit_buffer_0[335] = 8'h00;
    transmit_buffer_0[336] = 8'h00;
    transmit_buffer_0[337] = 8'h00;
    transmit_buffer_0[338] = 8'h00;
    transmit_buffer_0[339] = 8'h00;
    transmit_buffer_0[340] = 8'h00;
    transmit_buffer_0[341] = 8'h00;
    transmit_buffer_0[342] = 8'h00;
    transmit_buffer_0[343] = 8'h00;
    transmit_buffer_0[344] = 8'h00;
    transmit_buffer_0[345] = 8'h00;
    transmit_buffer_0[346] = 8'h00;
    transmit_buffer_0[347] = 8'h00;
    transmit_buffer_0[348] = 8'h00;
    transmit_buffer_0[349] = 8'h00;
    transmit_buffer_0[350] = 8'h00;
    transmit_buffer_0[351] = 8'h00;
    transmit_buffer_0[352] = 8'h00;
    transmit_buffer_0[353] = 8'h00;
    transmit_buffer_0[354] = 8'h00;
    transmit_buffer_0[355] = 8'h00;
    transmit_buffer_0[356] = 8'h00;
    transmit_buffer_0[357] = 8'h00;
    transmit_buffer_0[358] = 8'h00;
    transmit_buffer_0[359] = 8'h00;
    transmit_buffer_0[360] = 8'h00;
    transmit_buffer_0[361] = 8'h00;
    transmit_buffer_0[362] = 8'h00;
    transmit_buffer_0[363] = 8'h00;
    transmit_buffer_0[364] = 8'h00;
    transmit_buffer_0[365] = 8'h00;
    transmit_buffer_0[366] = 8'h00;
    transmit_buffer_0[367] = 8'h00;
    transmit_buffer_0[368] = 8'h00;
    transmit_buffer_0[369] = 8'h00;
    transmit_buffer_0[370] = 8'h00;
    transmit_buffer_0[371] = 8'h00;
    transmit_buffer_0[372] = 8'h00;
    transmit_buffer_0[373] = 8'h00;
    transmit_buffer_0[374] = 8'h00;
    transmit_buffer_0[375] = 8'h00;
    transmit_buffer_0[376] = 8'h00;
    transmit_buffer_0[377] = 8'h00;
    transmit_buffer_0[378] = 8'h00;
    transmit_buffer_0[379] = 8'h00;
    transmit_buffer_0[380] = 8'h00;
    transmit_buffer_0[381] = 8'h00;
    transmit_buffer_0[382] = 8'h00;
    transmit_buffer_0[383] = 8'h00;
    transmit_buffer_0[384] = 8'h00;
    transmit_buffer_0[385] = 8'h00;
    transmit_buffer_0[386] = 8'h00;
    transmit_buffer_0[387] = 8'h00;
    transmit_buffer_0[388] = 8'h00;
    transmit_buffer_0[389] = 8'h00;
    transmit_buffer_0[390] = 8'h00;
    transmit_buffer_0[391] = 8'h00;
    transmit_buffer_0[392] = 8'h00;
    transmit_buffer_0[393] = 8'h00;
    transmit_buffer_0[394] = 8'h00;
    transmit_buffer_0[395] = 8'h00;
    transmit_buffer_0[396] = 8'h00;
    transmit_buffer_0[397] = 8'h00;
    transmit_buffer_0[398] = 8'h00;
    transmit_buffer_0[399] = 8'h00;
    transmit_buffer_0[400] = 8'h00;
    transmit_buffer_0[401] = 8'h00;
    transmit_buffer_0[402] = 8'h00;
    transmit_buffer_0[403] = 8'h00;
    transmit_buffer_0[404] = 8'h00;
    transmit_buffer_0[405] = 8'h00;
    transmit_buffer_0[406] = 8'h00;
    transmit_buffer_0[407] = 8'h00;
    transmit_buffer_0[408] = 8'h00;
    transmit_buffer_0[409] = 8'h00;
    transmit_buffer_0[410] = 8'h00;
    transmit_buffer_0[411] = 8'h00;
    transmit_buffer_0[412] = 8'h00;
    transmit_buffer_0[413] = 8'h00;
    transmit_buffer_0[414] = 8'h00;
    transmit_buffer_0[415] = 8'h00;
    transmit_buffer_0[416] = 8'h00;
    transmit_buffer_0[417] = 8'h00;
    transmit_buffer_0[418] = 8'h00;
    transmit_buffer_0[419] = 8'h00;
    transmit_buffer_0[420] = 8'h00;
    transmit_buffer_0[421] = 8'h00;
    transmit_buffer_0[422] = 8'h00;
    transmit_buffer_0[423] = 8'h00;
    transmit_buffer_0[424] = 8'h00;
    transmit_buffer_0[425] = 8'h00;
    transmit_buffer_0[426] = 8'h00;
    transmit_buffer_0[427] = 8'h00;
    transmit_buffer_0[428] = 8'h00;
    transmit_buffer_0[429] = 8'h00;
    transmit_buffer_0[430] = 8'h00;
    transmit_buffer_0[431] = 8'h00;
    transmit_buffer_0[432] = 8'h00;
    transmit_buffer_0[433] = 8'h00;
    transmit_buffer_0[434] = 8'h00;
    transmit_buffer_0[435] = 8'h00;
    transmit_buffer_0[436] = 8'h00;
    transmit_buffer_0[437] = 8'h00;
    transmit_buffer_0[438] = 8'h00;
    transmit_buffer_0[439] = 8'h00;
    transmit_buffer_0[440] = 8'h00;
    transmit_buffer_0[441] = 8'h00;
    transmit_buffer_0[442] = 8'h00;
    transmit_buffer_0[443] = 8'h00;
    transmit_buffer_0[444] = 8'h00;
    transmit_buffer_0[445] = 8'h00;
    transmit_buffer_0[446] = 8'h00;
    transmit_buffer_0[447] = 8'h00;
    transmit_buffer_0[448] = 8'h00;
    transmit_buffer_0[449] = 8'h00;
    transmit_buffer_0[450] = 8'h00;
    transmit_buffer_0[451] = 8'h00;
    transmit_buffer_0[452] = 8'h00;
    transmit_buffer_0[453] = 8'h00;
    transmit_buffer_0[454] = 8'h00;
    transmit_buffer_0[455] = 8'h00;
    transmit_buffer_0[456] = 8'h00;
    transmit_buffer_0[457] = 8'h00;
    transmit_buffer_0[458] = 8'h00;
    transmit_buffer_0[459] = 8'h00;
    transmit_buffer_0[460] = 8'h00;
    transmit_buffer_0[461] = 8'h00;
    transmit_buffer_0[462] = 8'h00;
    transmit_buffer_0[463] = 8'h00;
    transmit_buffer_0[464] = 8'h00;
    transmit_buffer_0[465] = 8'h00;
    transmit_buffer_0[466] = 8'h00;
    transmit_buffer_0[467] = 8'h00;
    transmit_buffer_0[468] = 8'h00;
    transmit_buffer_0[469] = 8'h00;
    transmit_buffer_0[470] = 8'h00;
    transmit_buffer_0[471] = 8'h00;
    transmit_buffer_0[472] = 8'h00;
    transmit_buffer_0[473] = 8'h00;
    transmit_buffer_0[474] = 8'h00;
    transmit_buffer_0[475] = 8'h00;
    transmit_buffer_0[476] = 8'h00;
    transmit_buffer_0[477] = 8'h00;
    transmit_buffer_0[478] = 8'h00;
    transmit_buffer_0[479] = 8'h00;
    transmit_buffer_0[480] = 8'h00;
    transmit_buffer_0[481] = 8'h00;
    transmit_buffer_0[482] = 8'h00;
    transmit_buffer_0[483] = 8'h00;
    transmit_buffer_0[484] = 8'h00;
    transmit_buffer_0[485] = 8'h00;
    transmit_buffer_0[486] = 8'h00;
    transmit_buffer_0[487] = 8'h00;
    transmit_buffer_0[488] = 8'h00;
    transmit_buffer_0[489] = 8'h00;
    transmit_buffer_0[490] = 8'h00;
    transmit_buffer_0[491] = 8'h00;
    transmit_buffer_0[492] = 8'h00;
    transmit_buffer_0[493] = 8'h00;
    transmit_buffer_0[494] = 8'h00;
    transmit_buffer_0[495] = 8'h00;
    transmit_buffer_0[496] = 8'h00;
    transmit_buffer_0[497] = 8'h00;
    transmit_buffer_0[498] = 8'h00;
    transmit_buffer_0[499] = 8'h00;
    transmit_buffer_0[500] = 8'h00;
    transmit_buffer_0[501] = 8'h00;
    transmit_buffer_0[502] = 8'h00;
    transmit_buffer_0[503] = 8'h00;
    transmit_buffer_0[504] = 8'h00;
    transmit_buffer_0[505] = 8'h00;
    transmit_buffer_0[506] = 8'h00;
    transmit_buffer_0[507] = 8'h00;
    transmit_buffer_0[508] = 8'h00;
    transmit_buffer_0[509] = 8'h00;
    transmit_buffer_0[510] = 8'h00;
    transmit_buffer_0[511] = 8'h00;
  end
  always @(posedge usb_clk) begin
    if (transmit_buffer_0_w_en)
      transmit_buffer_0[transmit_buffer_0_w_addr] <= transmit_buffer_0_w_data;
  end
  reg [8:0] _0_;
  always @(posedge usb_clk) begin
    _0_ <= transmit_buffer_0_r_addr;
  end
  assign transmit_buffer_0_r_data = transmit_buffer_0[_0_];
  reg [7:0] transmit_buffer_1 [511:0];
  initial begin
    transmit_buffer_1[0] = 8'h00;
    transmit_buffer_1[1] = 8'h00;
    transmit_buffer_1[2] = 8'h00;
    transmit_buffer_1[3] = 8'h00;
    transmit_buffer_1[4] = 8'h00;
    transmit_buffer_1[5] = 8'h00;
    transmit_buffer_1[6] = 8'h00;
    transmit_buffer_1[7] = 8'h00;
    transmit_buffer_1[8] = 8'h00;
    transmit_buffer_1[9] = 8'h00;
    transmit_buffer_1[10] = 8'h00;
    transmit_buffer_1[11] = 8'h00;
    transmit_buffer_1[12] = 8'h00;
    transmit_buffer_1[13] = 8'h00;
    transmit_buffer_1[14] = 8'h00;
    transmit_buffer_1[15] = 8'h00;
    transmit_buffer_1[16] = 8'h00;
    transmit_buffer_1[17] = 8'h00;
    transmit_buffer_1[18] = 8'h00;
    transmit_buffer_1[19] = 8'h00;
    transmit_buffer_1[20] = 8'h00;
    transmit_buffer_1[21] = 8'h00;
    transmit_buffer_1[22] = 8'h00;
    transmit_buffer_1[23] = 8'h00;
    transmit_buffer_1[24] = 8'h00;
    transmit_buffer_1[25] = 8'h00;
    transmit_buffer_1[26] = 8'h00;
    transmit_buffer_1[27] = 8'h00;
    transmit_buffer_1[28] = 8'h00;
    transmit_buffer_1[29] = 8'h00;
    transmit_buffer_1[30] = 8'h00;
    transmit_buffer_1[31] = 8'h00;
    transmit_buffer_1[32] = 8'h00;
    transmit_buffer_1[33] = 8'h00;
    transmit_buffer_1[34] = 8'h00;
    transmit_buffer_1[35] = 8'h00;
    transmit_buffer_1[36] = 8'h00;
    transmit_buffer_1[37] = 8'h00;
    transmit_buffer_1[38] = 8'h00;
    transmit_buffer_1[39] = 8'h00;
    transmit_buffer_1[40] = 8'h00;
    transmit_buffer_1[41] = 8'h00;
    transmit_buffer_1[42] = 8'h00;
    transmit_buffer_1[43] = 8'h00;
    transmit_buffer_1[44] = 8'h00;
    transmit_buffer_1[45] = 8'h00;
    transmit_buffer_1[46] = 8'h00;
    transmit_buffer_1[47] = 8'h00;
    transmit_buffer_1[48] = 8'h00;
    transmit_buffer_1[49] = 8'h00;
    transmit_buffer_1[50] = 8'h00;
    transmit_buffer_1[51] = 8'h00;
    transmit_buffer_1[52] = 8'h00;
    transmit_buffer_1[53] = 8'h00;
    transmit_buffer_1[54] = 8'h00;
    transmit_buffer_1[55] = 8'h00;
    transmit_buffer_1[56] = 8'h00;
    transmit_buffer_1[57] = 8'h00;
    transmit_buffer_1[58] = 8'h00;
    transmit_buffer_1[59] = 8'h00;
    transmit_buffer_1[60] = 8'h00;
    transmit_buffer_1[61] = 8'h00;
    transmit_buffer_1[62] = 8'h00;
    transmit_buffer_1[63] = 8'h00;
    transmit_buffer_1[64] = 8'h00;
    transmit_buffer_1[65] = 8'h00;
    transmit_buffer_1[66] = 8'h00;
    transmit_buffer_1[67] = 8'h00;
    transmit_buffer_1[68] = 8'h00;
    transmit_buffer_1[69] = 8'h00;
    transmit_buffer_1[70] = 8'h00;
    transmit_buffer_1[71] = 8'h00;
    transmit_buffer_1[72] = 8'h00;
    transmit_buffer_1[73] = 8'h00;
    transmit_buffer_1[74] = 8'h00;
    transmit_buffer_1[75] = 8'h00;
    transmit_buffer_1[76] = 8'h00;
    transmit_buffer_1[77] = 8'h00;
    transmit_buffer_1[78] = 8'h00;
    transmit_buffer_1[79] = 8'h00;
    transmit_buffer_1[80] = 8'h00;
    transmit_buffer_1[81] = 8'h00;
    transmit_buffer_1[82] = 8'h00;
    transmit_buffer_1[83] = 8'h00;
    transmit_buffer_1[84] = 8'h00;
    transmit_buffer_1[85] = 8'h00;
    transmit_buffer_1[86] = 8'h00;
    transmit_buffer_1[87] = 8'h00;
    transmit_buffer_1[88] = 8'h00;
    transmit_buffer_1[89] = 8'h00;
    transmit_buffer_1[90] = 8'h00;
    transmit_buffer_1[91] = 8'h00;
    transmit_buffer_1[92] = 8'h00;
    transmit_buffer_1[93] = 8'h00;
    transmit_buffer_1[94] = 8'h00;
    transmit_buffer_1[95] = 8'h00;
    transmit_buffer_1[96] = 8'h00;
    transmit_buffer_1[97] = 8'h00;
    transmit_buffer_1[98] = 8'h00;
    transmit_buffer_1[99] = 8'h00;
    transmit_buffer_1[100] = 8'h00;
    transmit_buffer_1[101] = 8'h00;
    transmit_buffer_1[102] = 8'h00;
    transmit_buffer_1[103] = 8'h00;
    transmit_buffer_1[104] = 8'h00;
    transmit_buffer_1[105] = 8'h00;
    transmit_buffer_1[106] = 8'h00;
    transmit_buffer_1[107] = 8'h00;
    transmit_buffer_1[108] = 8'h00;
    transmit_buffer_1[109] = 8'h00;
    transmit_buffer_1[110] = 8'h00;
    transmit_buffer_1[111] = 8'h00;
    transmit_buffer_1[112] = 8'h00;
    transmit_buffer_1[113] = 8'h00;
    transmit_buffer_1[114] = 8'h00;
    transmit_buffer_1[115] = 8'h00;
    transmit_buffer_1[116] = 8'h00;
    transmit_buffer_1[117] = 8'h00;
    transmit_buffer_1[118] = 8'h00;
    transmit_buffer_1[119] = 8'h00;
    transmit_buffer_1[120] = 8'h00;
    transmit_buffer_1[121] = 8'h00;
    transmit_buffer_1[122] = 8'h00;
    transmit_buffer_1[123] = 8'h00;
    transmit_buffer_1[124] = 8'h00;
    transmit_buffer_1[125] = 8'h00;
    transmit_buffer_1[126] = 8'h00;
    transmit_buffer_1[127] = 8'h00;
    transmit_buffer_1[128] = 8'h00;
    transmit_buffer_1[129] = 8'h00;
    transmit_buffer_1[130] = 8'h00;
    transmit_buffer_1[131] = 8'h00;
    transmit_buffer_1[132] = 8'h00;
    transmit_buffer_1[133] = 8'h00;
    transmit_buffer_1[134] = 8'h00;
    transmit_buffer_1[135] = 8'h00;
    transmit_buffer_1[136] = 8'h00;
    transmit_buffer_1[137] = 8'h00;
    transmit_buffer_1[138] = 8'h00;
    transmit_buffer_1[139] = 8'h00;
    transmit_buffer_1[140] = 8'h00;
    transmit_buffer_1[141] = 8'h00;
    transmit_buffer_1[142] = 8'h00;
    transmit_buffer_1[143] = 8'h00;
    transmit_buffer_1[144] = 8'h00;
    transmit_buffer_1[145] = 8'h00;
    transmit_buffer_1[146] = 8'h00;
    transmit_buffer_1[147] = 8'h00;
    transmit_buffer_1[148] = 8'h00;
    transmit_buffer_1[149] = 8'h00;
    transmit_buffer_1[150] = 8'h00;
    transmit_buffer_1[151] = 8'h00;
    transmit_buffer_1[152] = 8'h00;
    transmit_buffer_1[153] = 8'h00;
    transmit_buffer_1[154] = 8'h00;
    transmit_buffer_1[155] = 8'h00;
    transmit_buffer_1[156] = 8'h00;
    transmit_buffer_1[157] = 8'h00;
    transmit_buffer_1[158] = 8'h00;
    transmit_buffer_1[159] = 8'h00;
    transmit_buffer_1[160] = 8'h00;
    transmit_buffer_1[161] = 8'h00;
    transmit_buffer_1[162] = 8'h00;
    transmit_buffer_1[163] = 8'h00;
    transmit_buffer_1[164] = 8'h00;
    transmit_buffer_1[165] = 8'h00;
    transmit_buffer_1[166] = 8'h00;
    transmit_buffer_1[167] = 8'h00;
    transmit_buffer_1[168] = 8'h00;
    transmit_buffer_1[169] = 8'h00;
    transmit_buffer_1[170] = 8'h00;
    transmit_buffer_1[171] = 8'h00;
    transmit_buffer_1[172] = 8'h00;
    transmit_buffer_1[173] = 8'h00;
    transmit_buffer_1[174] = 8'h00;
    transmit_buffer_1[175] = 8'h00;
    transmit_buffer_1[176] = 8'h00;
    transmit_buffer_1[177] = 8'h00;
    transmit_buffer_1[178] = 8'h00;
    transmit_buffer_1[179] = 8'h00;
    transmit_buffer_1[180] = 8'h00;
    transmit_buffer_1[181] = 8'h00;
    transmit_buffer_1[182] = 8'h00;
    transmit_buffer_1[183] = 8'h00;
    transmit_buffer_1[184] = 8'h00;
    transmit_buffer_1[185] = 8'h00;
    transmit_buffer_1[186] = 8'h00;
    transmit_buffer_1[187] = 8'h00;
    transmit_buffer_1[188] = 8'h00;
    transmit_buffer_1[189] = 8'h00;
    transmit_buffer_1[190] = 8'h00;
    transmit_buffer_1[191] = 8'h00;
    transmit_buffer_1[192] = 8'h00;
    transmit_buffer_1[193] = 8'h00;
    transmit_buffer_1[194] = 8'h00;
    transmit_buffer_1[195] = 8'h00;
    transmit_buffer_1[196] = 8'h00;
    transmit_buffer_1[197] = 8'h00;
    transmit_buffer_1[198] = 8'h00;
    transmit_buffer_1[199] = 8'h00;
    transmit_buffer_1[200] = 8'h00;
    transmit_buffer_1[201] = 8'h00;
    transmit_buffer_1[202] = 8'h00;
    transmit_buffer_1[203] = 8'h00;
    transmit_buffer_1[204] = 8'h00;
    transmit_buffer_1[205] = 8'h00;
    transmit_buffer_1[206] = 8'h00;
    transmit_buffer_1[207] = 8'h00;
    transmit_buffer_1[208] = 8'h00;
    transmit_buffer_1[209] = 8'h00;
    transmit_buffer_1[210] = 8'h00;
    transmit_buffer_1[211] = 8'h00;
    transmit_buffer_1[212] = 8'h00;
    transmit_buffer_1[213] = 8'h00;
    transmit_buffer_1[214] = 8'h00;
    transmit_buffer_1[215] = 8'h00;
    transmit_buffer_1[216] = 8'h00;
    transmit_buffer_1[217] = 8'h00;
    transmit_buffer_1[218] = 8'h00;
    transmit_buffer_1[219] = 8'h00;
    transmit_buffer_1[220] = 8'h00;
    transmit_buffer_1[221] = 8'h00;
    transmit_buffer_1[222] = 8'h00;
    transmit_buffer_1[223] = 8'h00;
    transmit_buffer_1[224] = 8'h00;
    transmit_buffer_1[225] = 8'h00;
    transmit_buffer_1[226] = 8'h00;
    transmit_buffer_1[227] = 8'h00;
    transmit_buffer_1[228] = 8'h00;
    transmit_buffer_1[229] = 8'h00;
    transmit_buffer_1[230] = 8'h00;
    transmit_buffer_1[231] = 8'h00;
    transmit_buffer_1[232] = 8'h00;
    transmit_buffer_1[233] = 8'h00;
    transmit_buffer_1[234] = 8'h00;
    transmit_buffer_1[235] = 8'h00;
    transmit_buffer_1[236] = 8'h00;
    transmit_buffer_1[237] = 8'h00;
    transmit_buffer_1[238] = 8'h00;
    transmit_buffer_1[239] = 8'h00;
    transmit_buffer_1[240] = 8'h00;
    transmit_buffer_1[241] = 8'h00;
    transmit_buffer_1[242] = 8'h00;
    transmit_buffer_1[243] = 8'h00;
    transmit_buffer_1[244] = 8'h00;
    transmit_buffer_1[245] = 8'h00;
    transmit_buffer_1[246] = 8'h00;
    transmit_buffer_1[247] = 8'h00;
    transmit_buffer_1[248] = 8'h00;
    transmit_buffer_1[249] = 8'h00;
    transmit_buffer_1[250] = 8'h00;
    transmit_buffer_1[251] = 8'h00;
    transmit_buffer_1[252] = 8'h00;
    transmit_buffer_1[253] = 8'h00;
    transmit_buffer_1[254] = 8'h00;
    transmit_buffer_1[255] = 8'h00;
    transmit_buffer_1[256] = 8'h00;
    transmit_buffer_1[257] = 8'h00;
    transmit_buffer_1[258] = 8'h00;
    transmit_buffer_1[259] = 8'h00;
    transmit_buffer_1[260] = 8'h00;
    transmit_buffer_1[261] = 8'h00;
    transmit_buffer_1[262] = 8'h00;
    transmit_buffer_1[263] = 8'h00;
    transmit_buffer_1[264] = 8'h00;
    transmit_buffer_1[265] = 8'h00;
    transmit_buffer_1[266] = 8'h00;
    transmit_buffer_1[267] = 8'h00;
    transmit_buffer_1[268] = 8'h00;
    transmit_buffer_1[269] = 8'h00;
    transmit_buffer_1[270] = 8'h00;
    transmit_buffer_1[271] = 8'h00;
    transmit_buffer_1[272] = 8'h00;
    transmit_buffer_1[273] = 8'h00;
    transmit_buffer_1[274] = 8'h00;
    transmit_buffer_1[275] = 8'h00;
    transmit_buffer_1[276] = 8'h00;
    transmit_buffer_1[277] = 8'h00;
    transmit_buffer_1[278] = 8'h00;
    transmit_buffer_1[279] = 8'h00;
    transmit_buffer_1[280] = 8'h00;
    transmit_buffer_1[281] = 8'h00;
    transmit_buffer_1[282] = 8'h00;
    transmit_buffer_1[283] = 8'h00;
    transmit_buffer_1[284] = 8'h00;
    transmit_buffer_1[285] = 8'h00;
    transmit_buffer_1[286] = 8'h00;
    transmit_buffer_1[287] = 8'h00;
    transmit_buffer_1[288] = 8'h00;
    transmit_buffer_1[289] = 8'h00;
    transmit_buffer_1[290] = 8'h00;
    transmit_buffer_1[291] = 8'h00;
    transmit_buffer_1[292] = 8'h00;
    transmit_buffer_1[293] = 8'h00;
    transmit_buffer_1[294] = 8'h00;
    transmit_buffer_1[295] = 8'h00;
    transmit_buffer_1[296] = 8'h00;
    transmit_buffer_1[297] = 8'h00;
    transmit_buffer_1[298] = 8'h00;
    transmit_buffer_1[299] = 8'h00;
    transmit_buffer_1[300] = 8'h00;
    transmit_buffer_1[301] = 8'h00;
    transmit_buffer_1[302] = 8'h00;
    transmit_buffer_1[303] = 8'h00;
    transmit_buffer_1[304] = 8'h00;
    transmit_buffer_1[305] = 8'h00;
    transmit_buffer_1[306] = 8'h00;
    transmit_buffer_1[307] = 8'h00;
    transmit_buffer_1[308] = 8'h00;
    transmit_buffer_1[309] = 8'h00;
    transmit_buffer_1[310] = 8'h00;
    transmit_buffer_1[311] = 8'h00;
    transmit_buffer_1[312] = 8'h00;
    transmit_buffer_1[313] = 8'h00;
    transmit_buffer_1[314] = 8'h00;
    transmit_buffer_1[315] = 8'h00;
    transmit_buffer_1[316] = 8'h00;
    transmit_buffer_1[317] = 8'h00;
    transmit_buffer_1[318] = 8'h00;
    transmit_buffer_1[319] = 8'h00;
    transmit_buffer_1[320] = 8'h00;
    transmit_buffer_1[321] = 8'h00;
    transmit_buffer_1[322] = 8'h00;
    transmit_buffer_1[323] = 8'h00;
    transmit_buffer_1[324] = 8'h00;
    transmit_buffer_1[325] = 8'h00;
    transmit_buffer_1[326] = 8'h00;
    transmit_buffer_1[327] = 8'h00;
    transmit_buffer_1[328] = 8'h00;
    transmit_buffer_1[329] = 8'h00;
    transmit_buffer_1[330] = 8'h00;
    transmit_buffer_1[331] = 8'h00;
    transmit_buffer_1[332] = 8'h00;
    transmit_buffer_1[333] = 8'h00;
    transmit_buffer_1[334] = 8'h00;
    transmit_buffer_1[335] = 8'h00;
    transmit_buffer_1[336] = 8'h00;
    transmit_buffer_1[337] = 8'h00;
    transmit_buffer_1[338] = 8'h00;
    transmit_buffer_1[339] = 8'h00;
    transmit_buffer_1[340] = 8'h00;
    transmit_buffer_1[341] = 8'h00;
    transmit_buffer_1[342] = 8'h00;
    transmit_buffer_1[343] = 8'h00;
    transmit_buffer_1[344] = 8'h00;
    transmit_buffer_1[345] = 8'h00;
    transmit_buffer_1[346] = 8'h00;
    transmit_buffer_1[347] = 8'h00;
    transmit_buffer_1[348] = 8'h00;
    transmit_buffer_1[349] = 8'h00;
    transmit_buffer_1[350] = 8'h00;
    transmit_buffer_1[351] = 8'h00;
    transmit_buffer_1[352] = 8'h00;
    transmit_buffer_1[353] = 8'h00;
    transmit_buffer_1[354] = 8'h00;
    transmit_buffer_1[355] = 8'h00;
    transmit_buffer_1[356] = 8'h00;
    transmit_buffer_1[357] = 8'h00;
    transmit_buffer_1[358] = 8'h00;
    transmit_buffer_1[359] = 8'h00;
    transmit_buffer_1[360] = 8'h00;
    transmit_buffer_1[361] = 8'h00;
    transmit_buffer_1[362] = 8'h00;
    transmit_buffer_1[363] = 8'h00;
    transmit_buffer_1[364] = 8'h00;
    transmit_buffer_1[365] = 8'h00;
    transmit_buffer_1[366] = 8'h00;
    transmit_buffer_1[367] = 8'h00;
    transmit_buffer_1[368] = 8'h00;
    transmit_buffer_1[369] = 8'h00;
    transmit_buffer_1[370] = 8'h00;
    transmit_buffer_1[371] = 8'h00;
    transmit_buffer_1[372] = 8'h00;
    transmit_buffer_1[373] = 8'h00;
    transmit_buffer_1[374] = 8'h00;
    transmit_buffer_1[375] = 8'h00;
    transmit_buffer_1[376] = 8'h00;
    transmit_buffer_1[377] = 8'h00;
    transmit_buffer_1[378] = 8'h00;
    transmit_buffer_1[379] = 8'h00;
    transmit_buffer_1[380] = 8'h00;
    transmit_buffer_1[381] = 8'h00;
    transmit_buffer_1[382] = 8'h00;
    transmit_buffer_1[383] = 8'h00;
    transmit_buffer_1[384] = 8'h00;
    transmit_buffer_1[385] = 8'h00;
    transmit_buffer_1[386] = 8'h00;
    transmit_buffer_1[387] = 8'h00;
    transmit_buffer_1[388] = 8'h00;
    transmit_buffer_1[389] = 8'h00;
    transmit_buffer_1[390] = 8'h00;
    transmit_buffer_1[391] = 8'h00;
    transmit_buffer_1[392] = 8'h00;
    transmit_buffer_1[393] = 8'h00;
    transmit_buffer_1[394] = 8'h00;
    transmit_buffer_1[395] = 8'h00;
    transmit_buffer_1[396] = 8'h00;
    transmit_buffer_1[397] = 8'h00;
    transmit_buffer_1[398] = 8'h00;
    transmit_buffer_1[399] = 8'h00;
    transmit_buffer_1[400] = 8'h00;
    transmit_buffer_1[401] = 8'h00;
    transmit_buffer_1[402] = 8'h00;
    transmit_buffer_1[403] = 8'h00;
    transmit_buffer_1[404] = 8'h00;
    transmit_buffer_1[405] = 8'h00;
    transmit_buffer_1[406] = 8'h00;
    transmit_buffer_1[407] = 8'h00;
    transmit_buffer_1[408] = 8'h00;
    transmit_buffer_1[409] = 8'h00;
    transmit_buffer_1[410] = 8'h00;
    transmit_buffer_1[411] = 8'h00;
    transmit_buffer_1[412] = 8'h00;
    transmit_buffer_1[413] = 8'h00;
    transmit_buffer_1[414] = 8'h00;
    transmit_buffer_1[415] = 8'h00;
    transmit_buffer_1[416] = 8'h00;
    transmit_buffer_1[417] = 8'h00;
    transmit_buffer_1[418] = 8'h00;
    transmit_buffer_1[419] = 8'h00;
    transmit_buffer_1[420] = 8'h00;
    transmit_buffer_1[421] = 8'h00;
    transmit_buffer_1[422] = 8'h00;
    transmit_buffer_1[423] = 8'h00;
    transmit_buffer_1[424] = 8'h00;
    transmit_buffer_1[425] = 8'h00;
    transmit_buffer_1[426] = 8'h00;
    transmit_buffer_1[427] = 8'h00;
    transmit_buffer_1[428] = 8'h00;
    transmit_buffer_1[429] = 8'h00;
    transmit_buffer_1[430] = 8'h00;
    transmit_buffer_1[431] = 8'h00;
    transmit_buffer_1[432] = 8'h00;
    transmit_buffer_1[433] = 8'h00;
    transmit_buffer_1[434] = 8'h00;
    transmit_buffer_1[435] = 8'h00;
    transmit_buffer_1[436] = 8'h00;
    transmit_buffer_1[437] = 8'h00;
    transmit_buffer_1[438] = 8'h00;
    transmit_buffer_1[439] = 8'h00;
    transmit_buffer_1[440] = 8'h00;
    transmit_buffer_1[441] = 8'h00;
    transmit_buffer_1[442] = 8'h00;
    transmit_buffer_1[443] = 8'h00;
    transmit_buffer_1[444] = 8'h00;
    transmit_buffer_1[445] = 8'h00;
    transmit_buffer_1[446] = 8'h00;
    transmit_buffer_1[447] = 8'h00;
    transmit_buffer_1[448] = 8'h00;
    transmit_buffer_1[449] = 8'h00;
    transmit_buffer_1[450] = 8'h00;
    transmit_buffer_1[451] = 8'h00;
    transmit_buffer_1[452] = 8'h00;
    transmit_buffer_1[453] = 8'h00;
    transmit_buffer_1[454] = 8'h00;
    transmit_buffer_1[455] = 8'h00;
    transmit_buffer_1[456] = 8'h00;
    transmit_buffer_1[457] = 8'h00;
    transmit_buffer_1[458] = 8'h00;
    transmit_buffer_1[459] = 8'h00;
    transmit_buffer_1[460] = 8'h00;
    transmit_buffer_1[461] = 8'h00;
    transmit_buffer_1[462] = 8'h00;
    transmit_buffer_1[463] = 8'h00;
    transmit_buffer_1[464] = 8'h00;
    transmit_buffer_1[465] = 8'h00;
    transmit_buffer_1[466] = 8'h00;
    transmit_buffer_1[467] = 8'h00;
    transmit_buffer_1[468] = 8'h00;
    transmit_buffer_1[469] = 8'h00;
    transmit_buffer_1[470] = 8'h00;
    transmit_buffer_1[471] = 8'h00;
    transmit_buffer_1[472] = 8'h00;
    transmit_buffer_1[473] = 8'h00;
    transmit_buffer_1[474] = 8'h00;
    transmit_buffer_1[475] = 8'h00;
    transmit_buffer_1[476] = 8'h00;
    transmit_buffer_1[477] = 8'h00;
    transmit_buffer_1[478] = 8'h00;
    transmit_buffer_1[479] = 8'h00;
    transmit_buffer_1[480] = 8'h00;
    transmit_buffer_1[481] = 8'h00;
    transmit_buffer_1[482] = 8'h00;
    transmit_buffer_1[483] = 8'h00;
    transmit_buffer_1[484] = 8'h00;
    transmit_buffer_1[485] = 8'h00;
    transmit_buffer_1[486] = 8'h00;
    transmit_buffer_1[487] = 8'h00;
    transmit_buffer_1[488] = 8'h00;
    transmit_buffer_1[489] = 8'h00;
    transmit_buffer_1[490] = 8'h00;
    transmit_buffer_1[491] = 8'h00;
    transmit_buffer_1[492] = 8'h00;
    transmit_buffer_1[493] = 8'h00;
    transmit_buffer_1[494] = 8'h00;
    transmit_buffer_1[495] = 8'h00;
    transmit_buffer_1[496] = 8'h00;
    transmit_buffer_1[497] = 8'h00;
    transmit_buffer_1[498] = 8'h00;
    transmit_buffer_1[499] = 8'h00;
    transmit_buffer_1[500] = 8'h00;
    transmit_buffer_1[501] = 8'h00;
    transmit_buffer_1[502] = 8'h00;
    transmit_buffer_1[503] = 8'h00;
    transmit_buffer_1[504] = 8'h00;
    transmit_buffer_1[505] = 8'h00;
    transmit_buffer_1[506] = 8'h00;
    transmit_buffer_1[507] = 8'h00;
    transmit_buffer_1[508] = 8'h00;
    transmit_buffer_1[509] = 8'h00;
    transmit_buffer_1[510] = 8'h00;
    transmit_buffer_1[511] = 8'h00;
  end
  always @(posedge usb_clk) begin
    if (transmit_buffer_1_w_en)
      transmit_buffer_1[transmit_buffer_1_w_addr] <= transmit_buffer_1_w_data;
  end
  reg [8:0] _1_;
  always @(posedge usb_clk) begin
    _1_ <= transmit_buffer_1_r_addr;
  end
  assign transmit_buffer_1_r_data = transmit_buffer_1[_1_];
  assign \$100  = generate_zlps &  \$98 ;
  assign \$102  = \$100  &  stream_ended_in_buffer1;
  assign \$104  = ~  ready;
  assign \$106  = \$signal$27  ==  10'h200;
  assign \$108  = generate_zlps &  \$106 ;
  assign \$110  = \$108  &  stream_ended_in_buffer1;
  assign \$112  = ~  ready;
  assign \$114  = \$signal  +  1'h1;
  assign \$116  = \$114  ==  10'h200;
  assign \$118  = \$116  |  last;
  assign \$11  = \$signal  +  1'h1;
  assign \$120  = valid &  \$118 ;
  assign \$122  = \$112  |  \$120 ;
  assign \$124  = ~  data_pid[0];
  assign \$126  = ~  data_pid[0];
  assign \$128  = \$signal$27  ==  10'h200;
  assign \$130  = generate_zlps &  \$128 ;
  assign \$132  = \$130  &  stream_ended_in_buffer1;
  assign \$134  = ~  ready;
  assign \$136  = \$signal$27  +  1'h1;
  assign \$138  = \$136  ==  10'h200;
  assign \$13  = \$11  ==  10'h200;
  assign \$140  = \$138  |  last;
  assign \$142  = valid &  \$140 ;
  assign \$144  = \$134  |  \$142 ;
  assign \$146  = ~  data_pid[0];
  assign \$148  = ~  data_pid[0];
  assign \$156  = ~  buffer_toggle;
  assign \$15  = \$13  |  last;
  assign \$159  = send_position +  1'h1;
  assign \$161  = ~  buffer_toggle;
  assign \$164  = send_position +  1'h1;
  assign \$167  = send_position +  1'h1;
  assign \$169  = ~  buffer_toggle;
  assign \$171  = \$signal  !=  10'h200;
  assign \$173  = ~  stream_ended_in_buffer0;
  assign \$175  = \$171  &  \$173 ;
  assign \$177  = \$signal$27  !=  10'h200;
  assign \$17  = valid &  \$15 ;
  assign \$179  = ~  stream_ended_in_buffer1;
  assign \$181  = \$177  &  \$179 ;
  assign \$183  = valid &  ready;
  assign \$185  = valid &  ready;
  assign \$187  = valid &  ready;
  assign \$190  = \$signal  +  1'h1;
  assign \$193  = \$signal$27  +  1'h1;
  assign \$195  = ~  buffer_toggle;
  assign \$197  = last &  transmit_buffer_0_w_en;
  assign \$19  = \$signal  +  1'h1;
  assign \$199  = last &  transmit_buffer_1_w_en;
  assign \$201  = \$signal  +  1'h1;
  assign \$203  = \$201  ==  10'h200;
  assign \$205  = \$203  |  last;
  assign \$207  = valid &  \$205 ;
  assign \$209  = \$signal  +  1'h1;
  assign \$211  = \$209  ==  10'h200;
  assign \$213  = \$211  |  last;
  assign \$217  = \$signal$27  +  1'h1;
  assign \$21  = \$19  ==  10'h200;
  assign \$219  = \$217  ==  10'h200;
  assign \$221  = \$219  |  last;
  assign \$223  = valid &  \$221 ;
  assign \$225  = \$signal$27  +  1'h1;
  assign \$227  = \$225  ==  10'h200;
  assign \$229  = \$227  |  last;
  assign \$233  = active &  is_in;
  assign \$235  = \$233  &  ready_for_response;
  assign \$238  = ~  buffer_toggle;
  assign \$23  = \$21  |  last;
  assign \$240  = |  \$signal ;
  assign \$242  = |  \$signal$27 ;
  assign \$244  = ~  buffer_toggle;
  assign \$246  = \$signal  ==  10'h200;
  assign \$248  = generate_zlps &  \$246 ;
  assign \$250  = \$248  &  stream_ended_in_buffer0;
  assign \$252  = ~  ready;
  assign \$254  = \$signal  ==  10'h200;
  assign \$256  = generate_zlps &  \$254 ;
  assign \$258  = \$256  &  stream_ended_in_buffer0;
  assign \$25  = ~  data_pid[0];
  assign \$260  = ~  ready;
  assign \$262  = \$signal  +  1'h1;
  assign \$264  = \$262  ==  10'h200;
  assign \$266  = \$264  |  last;
  assign \$268  = valid &  \$266 ;
  assign \$270  = \$260  |  \$268 ;
  assign \$272  = \$signal  ==  10'h200;
  assign \$274  = generate_zlps &  \$272 ;
  assign \$276  = \$274  &  stream_ended_in_buffer0;
  assign \$278  = ~  ready;
  assign \$280  = \$signal$27  +  1'h1;
  assign \$282  = \$280  ==  10'h200;
  assign \$284  = \$282  |  last;
  assign \$286  = valid &  \$284 ;
  assign \$288  = \$278  |  \$286 ;
  assign \$28  = \$signal$27  +  1'h1;
  assign \$290  = \$signal$27  ==  10'h200;
  assign \$292  = generate_zlps &  \$290 ;
  assign \$294  = \$292  &  stream_ended_in_buffer1;
  assign \$296  = ~  ready;
  assign \$298  = \$signal$27  ==  10'h200;
  assign \$300  = generate_zlps &  \$298 ;
  assign \$302  = \$300  &  stream_ended_in_buffer1;
  assign \$304  = ~  ready;
  assign \$306  = \$signal  +  1'h1;
  assign \$308  = \$306  ==  10'h200;
  assign \$30  = \$28  ==  10'h200;
  assign \$310  = \$308  |  last;
  assign \$312  = valid &  \$310 ;
  assign \$314  = \$304  |  \$312 ;
  assign \$316  = \$signal$27  ==  10'h200;
  assign \$318  = generate_zlps &  \$316 ;
  assign \$320  = \$318  &  stream_ended_in_buffer1;
  assign \$322  = ~  ready;
  assign \$324  = \$signal$27  +  1'h1;
  assign \$326  = \$324  ==  10'h200;
  assign \$328  = \$326  |  last;
  assign \$32  = \$30  |  last;
  assign \$330  = valid &  \$328 ;
  assign \$332  = \$322  |  \$330 ;
  assign \$334  = active &  is_in;
  assign \$336  = \$334  &  ready_for_response;
  assign \$338  = \$signal  +  1'h1;
  assign \$340  = \$338  ==  10'h200;
  assign \$342  = \$340  |  last;
  assign \$344  = valid &  \$342 ;
  assign \$346  = \$signal  +  1'h1;
  assign \$348  = \$346  ==  10'h200;
  assign \$34  = valid &  \$32 ;
  assign \$350  = \$348  |  last;
  assign \$352  = \$signal$27  +  1'h1;
  assign \$354  = \$352  ==  10'h200;
  assign \$356  = \$354  |  last;
  assign \$358  = valid &  \$356 ;
  assign \$360  = \$signal$27  +  1'h1;
  assign \$362  = \$360  ==  10'h200;
  assign \$364  = \$362  |  last;
  assign \$366  = active &  is_in;
  assign \$368  = \$366  &  ready_for_response;
  assign \$36  = \$signal$27  +  1'h1;
  assign \$371  = ~  buffer_toggle;
  assign \$373  = |  \$signal ;
  assign \$375  = |  \$signal$27 ;
  assign \$377  = send_position +  1'h1;
  assign \$379  = ~  buffer_toggle;
  assign \$381  = send_position +  1'h1;
  assign \$383  = \$381  ==  \$signal ;
  assign \$385  = send_position +  1'h1;
  assign \$387  = \$385  ==  \$signal$27 ;
  assign \$38  = \$36  ==  10'h200;
  assign \$389  = ~  buffer_toggle;
  assign \$391  = \$signal  ==  10'h200;
  assign \$393  = generate_zlps &  \$391 ;
  assign \$395  = \$393  &  stream_ended_in_buffer0;
  assign \$397  = ~  ready;
  assign \$399  = \$signal  ==  10'h200;
  assign \$401  = generate_zlps &  \$399 ;
  assign \$403  = \$401  &  stream_ended_in_buffer0;
  assign \$405  = ~  ready;
  assign \$407  = \$signal  +  1'h1;
  assign \$40  = \$38  |  last;
  assign \$409  = \$407  ==  10'h200;
  assign \$411  = \$409  |  last;
  assign \$413  = valid &  \$411 ;
  assign \$415  = \$405  |  \$413 ;
  assign \$417  = \$signal  ==  10'h200;
  assign \$419  = generate_zlps &  \$417 ;
  assign \$421  = \$419  &  stream_ended_in_buffer0;
  assign \$423  = ~  ready;
  assign \$425  = \$signal$27  +  1'h1;
  assign \$427  = \$425  ==  10'h200;
  assign \$42  = ~  data_pid[0];
  assign \$429  = \$427  |  last;
  assign \$431  = valid &  \$429 ;
  assign \$433  = \$423  |  \$431 ;
  assign \$435  = \$signal$27  ==  10'h200;
  assign \$437  = generate_zlps &  \$435 ;
  assign \$439  = \$437  &  stream_ended_in_buffer1;
  assign \$441  = ~  ready;
  assign \$443  = \$signal$27  ==  10'h200;
  assign \$445  = generate_zlps &  \$443 ;
  assign \$447  = \$445  &  stream_ended_in_buffer1;
  assign \$44  = ~  buffer_toggle;
  assign \$449  = ~  ready;
  assign \$451  = \$signal  +  1'h1;
  assign \$453  = \$451  ==  10'h200;
  assign \$455  = \$453  |  last;
  assign \$457  = valid &  \$455 ;
  assign \$459  = \$449  |  \$457 ;
  assign \$461  = \$signal$27  ==  10'h200;
  assign \$463  = generate_zlps &  \$461 ;
  assign \$465  = \$463  &  stream_ended_in_buffer1;
  assign \$467  = ~  ready;
  assign \$46  = \$signal  ==  10'h200;
  assign \$469  = \$signal$27  +  1'h1;
  assign \$471  = \$469  ==  10'h200;
  assign \$473  = \$471  |  last;
  assign \$475  = valid &  \$473 ;
  assign \$477  = \$467  |  \$475 ;
  assign \$479  = \$signal  +  1'h1;
  assign \$481  = \$479  ==  10'h200;
  assign \$483  = \$481  |  last;
  assign \$485  = valid &  \$483 ;
  assign \$487  = \$signal  +  1'h1;
  assign \$48  = generate_zlps &  \$46 ;
  assign \$489  = \$487  ==  10'h200;
  assign \$491  = \$489  |  last;
  assign \$495  = \$signal$27  +  1'h1;
  assign \$497  = \$495  ==  10'h200;
  assign \$499  = \$497  |  last;
  assign \$501  = valid &  \$499 ;
  assign \$503  = \$signal$27  +  1'h1;
  assign \$505  = \$503  ==  10'h200;
  assign \$507  = \$505  |  last;
  assign \$50  = \$48  &  stream_ended_in_buffer0;
  assign \$511  = ~  buffer_toggle;
  assign \$513  = \$signal  ==  10'h200;
  assign \$515  = generate_zlps &  \$513 ;
  assign \$517  = \$515  &  stream_ended_in_buffer0;
  assign \$519  = ~  ready;
  assign \$521  = \$signal  ==  10'h200;
  assign \$523  = generate_zlps &  \$521 ;
  assign \$525  = \$523  &  stream_ended_in_buffer0;
  assign \$527  = ~  ready;
  assign \$52  = ~  ready;
  assign \$529  = \$signal  +  1'h1;
  assign \$531  = \$529  ==  10'h200;
  assign \$533  = \$531  |  last;
  assign \$535  = valid &  \$533 ;
  assign \$537  = \$527  |  \$535 ;
  assign \$539  = \$signal  ==  10'h200;
  assign \$541  = generate_zlps &  \$539 ;
  assign \$543  = \$541  &  stream_ended_in_buffer0;
  assign \$545  = ~  ready;
  assign \$547  = \$signal$27  +  1'h1;
  assign \$54  = \$signal  ==  10'h200;
  assign \$549  = \$547  ==  10'h200;
  assign \$551  = \$549  |  last;
  assign \$553  = valid &  \$551 ;
  assign \$555  = \$545  |  \$553 ;
  assign \$557  = \$signal$27  ==  10'h200;
  assign \$559  = generate_zlps &  \$557 ;
  assign \$561  = \$559  &  stream_ended_in_buffer1;
  assign \$563  = ~  ready;
  assign \$565  = \$signal$27  ==  10'h200;
  assign \$567  = generate_zlps &  \$565 ;
  assign \$56  = generate_zlps &  \$54 ;
  assign \$569  = \$567  &  stream_ended_in_buffer1;
  assign \$571  = ~  ready;
  assign \$573  = \$signal  +  1'h1;
  assign \$575  = \$573  ==  10'h200;
  assign \$577  = \$575  |  last;
  assign \$579  = valid &  \$577 ;
  assign \$581  = \$571  |  \$579 ;
  assign \$583  = \$signal$27  ==  10'h200;
  assign \$585  = generate_zlps &  \$583 ;
  assign \$587  = \$585  &  stream_ended_in_buffer1;
  assign \$58  = \$56  &  stream_ended_in_buffer0;
  assign \$589  = ~  ready;
  assign \$591  = \$signal$27  +  1'h1;
  assign \$593  = \$591  ==  10'h200;
  assign \$595  = \$593  |  last;
  assign \$597  = valid &  \$595 ;
  assign \$599  = \$589  |  \$597 ;
  assign \$602  = send_position +  1'h1;
  assign \$604  = active &  is_in;
  assign \$606  = \$604  &  ready_for_response;
  assign \$60  = ~  ready;
  assign \$609  = ~  buffer_toggle;
  assign \$611  = |  \$signal ;
  assign \$613  = |  \$signal$27 ;
  assign \$615  = active &  is_in;
  assign \$617  = \$615  &  ready_for_response;
  assign \$620  = ~  buffer_toggle;
  assign \$622  = |  \$signal ;
  assign \$624  = |  \$signal$27 ;
  assign \$626  = active &  is_in;
  assign \$628  = \$626  &  ready_for_response;
  assign \$62  = \$signal  +  1'h1;
  assign \$631  = ~  buffer_toggle;
  assign \$633  = |  \$signal ;
  assign \$635  = |  \$signal$27 ;
  assign \$637  = send_position +  1'h1;
  assign \$639  = ~  buffer_toggle;
  assign \$641  = send_position +  1'h1;
  assign \$643  = \$641  ==  \$signal ;
  assign \$645  = send_position +  1'h1;
  assign \$647  = \$645  ==  \$signal$27 ;
  always @(posedge usb_clk)
    data_pid <= \data_pid$next ;
  assign \$64  = \$62  ==  10'h200;
  always @(posedge usb_clk)
    \$signal  <= \$signal$next ;
  always @(posedge usb_clk)
    \$signal$27  <= \$signal$27$next ;
  always @(posedge usb_clk)
    stream_ended_in_buffer0 <= \stream_ended_in_buffer0$next ;
  always @(posedge usb_clk)
    stream_ended_in_buffer1 <= \stream_ended_in_buffer1$next ;
  always @(posedge usb_clk)
    fsm_state <= \fsm_state$next ;
  always @(posedge usb_clk)
    buffer_toggle <= \buffer_toggle$next ;
  always @(posedge usb_clk)
    send_position <= \send_position$next ;
  always @(posedge usb_clk)
    first <= \first$next ;
  assign \$66  = \$64  |  last;
  assign \$68  = valid &  \$66 ;
  assign \$70  = \$60  |  \$68 ;
  assign \$72  = ~  data_pid[0];
  assign \$74  = ~  data_pid[0];
  assign \$76  = \$signal  ==  10'h200;
  assign \$78  = generate_zlps &  \$76 ;
  assign \$80  = \$78  &  stream_ended_in_buffer0;
  assign \$82  = ~  ready;
  assign \$84  = \$signal$27  +  1'h1;
  assign \$86  = \$84  ==  10'h200;
  assign \$88  = \$86  |  last;
  assign \$90  = valid &  \$88 ;
  assign \$92  = \$82  |  \$90 ;
  assign \$94  = ~  data_pid[0];
  assign \$96  = ~  data_pid[0];
  assign \$98  = \$signal$27  ==  10'h200;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$31 ) begin end
    \data_pid$next  = data_pid;
    casez (reset_sequence)
      1'h1:
          \data_pid$next  = \$7 ;
    endcase
    casez (fsm_state)
      2'h0:
          casez (buffer_toggle)
            1'h0:
                casez (\$17 )
                  1'h1:
                      casez (\$23 )
                        1'h1:
                            \data_pid$next [0] = \$25 ;
                      endcase
                endcase
            1'h?:
                casez (\$34 )
                  1'h1:
                      casez (\$40 )
                        1'h1:
                            \data_pid$next [0] = \$42 ;
                      endcase
                endcase
          endcase
      2'h1:
          ;
      2'h2:
          ;
      2'h3:
          casez (ack)
            1'h1:
                casez (\$44 )
                  1'h0:
                      casez (buffer_toggle)
                        1'h0:
                            casez ({ \$70 , \$58  })
                              2'b?1:
                                  \data_pid$next [0] = \$72 ;
                              2'b1?:
                                  \data_pid$next [0] = \$74 ;
                            endcase
                        1'h?:
                            casez ({ \$92 , \$80  })
                              2'b?1:
                                  \data_pid$next [0] = \$94 ;
                              2'b1?:
                                  \data_pid$next [0] = \$96 ;
                            endcase
                      endcase
                  1'h?:
                      casez (buffer_toggle)
                        1'h0:
                            casez ({ \$122 , \$110  })
                              2'b?1:
                                  \data_pid$next [0] = \$124 ;
                              2'b1?:
                                  \data_pid$next [0] = \$126 ;
                            endcase
                        1'h?:
                            casez ({ \$144 , \$132  })
                              2'b?1:
                                  \data_pid$next [0] = \$146 ;
                              2'b1?:
                                  \data_pid$next [0] = \$148 ;
                            endcase
                      endcase
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \data_pid$next  = 2'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$31 ) begin end
    \$signal$next  = \$signal ;
    \$signal$27$next  = \$signal$27 ;
    casez (buffer_toggle)
      1'h0:
          casez (transmit_buffer_0_w_en)
            1'h1:
                \$signal$next  = \$190 [9:0];
          endcase
      1'h?:
          casez (transmit_buffer_1_w_en)
            1'h1:
                \$signal$27$next  = \$193 [9:0];
          endcase
    endcase
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          ;
      2'h2:
          ;
      2'h3:
          casez (ack)
            1'h1:
                casez (\$195 )
                  1'h0:
                      \$signal$next  = 10'h000;
                  1'h?:
                      \$signal$27$next  = 10'h000;
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
        begin
          \$signal$next  = 10'h000;
          \$signal$27$next  = 10'h000;
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$31 ) begin end
    \stream_ended_in_buffer0$next  = stream_ended_in_buffer0;
    \stream_ended_in_buffer1$next  = stream_ended_in_buffer1;
    casez (buffer_toggle)
      1'h0:
          casez (\$197 )
            1'h1:
                \stream_ended_in_buffer0$next  = 1'h1;
          endcase
      1'h?:
          casez (\$199 )
            1'h1:
                \stream_ended_in_buffer1$next  = 1'h1;
          endcase
    endcase
    casez (fsm_state)
      2'h0:
          casez (buffer_toggle)
            1'h0:
                casez (\$207 )
                  1'h1:
                      casez (\$213 )
                        1'h1:
                            casez (\$215 )
                              1'h0:
                                  \stream_ended_in_buffer0$next  = 1'h0;
                              1'h?:
                                  \stream_ended_in_buffer1$next  = 1'h0;
                            endcase
                      endcase
                endcase
            1'h?:
                casez (\$223 )
                  1'h1:
                      casez (\$229 )
                        1'h1:
                            casez (\$231 )
                              1'h0:
                                  \stream_ended_in_buffer0$next  = 1'h0;
                              1'h?:
                                  \stream_ended_in_buffer1$next  = 1'h0;
                            endcase
                      endcase
                endcase
          endcase
      2'h1:
          casez (\$235 )
            1'h1:
                casez (\$238 )
                  1'h0:
                      casez (\$240 )
                        1'h1:
                            ;
                        default:
                            \stream_ended_in_buffer0$next  = 1'h0;
                      endcase
                  1'h?:
                      casez (\$242 )
                        1'h1:
                            ;
                        default:
                            \stream_ended_in_buffer1$next  = 1'h0;
                      endcase
                endcase
          endcase
      2'h2:
          ;
      2'h3:
          casez (ack)
            1'h1:
                casez (\$244 )
                  1'h0:
                      casez (buffer_toggle)
                        1'h0:
                            casez ({ \$270 , \$258  })
                              2'b?1:
                                  ;
                              2'b1?:
                                  \stream_ended_in_buffer0$next  = 1'h0;
                            endcase
                        1'h?:
                            casez ({ \$288 , \$276  })
                              2'b?1:
                                  ;
                              2'b1?:
                                  \stream_ended_in_buffer0$next  = 1'h0;
                            endcase
                      endcase
                  1'h?:
                      casez (buffer_toggle)
                        1'h0:
                            casez ({ \$314 , \$302  })
                              2'b?1:
                                  ;
                              2'b1?:
                                  \stream_ended_in_buffer1$next  = 1'h0;
                            endcase
                        1'h?:
                            casez ({ \$332 , \$320  })
                              2'b?1:
                                  ;
                              2'b1?:
                                  \stream_ended_in_buffer1$next  = 1'h0;
                            endcase
                      endcase
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
        begin
          \stream_ended_in_buffer0$next  = 1'h0;
          \stream_ended_in_buffer1$next  = 1'h0;
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$31 ) begin end
    nak = 1'h0;
    casez (fsm_state)
      2'h0:
          nak = \$336 ;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$31 ) begin end
    \fsm_state$next  = fsm_state;
    casez (fsm_state)
      2'h0:
          casez (buffer_toggle)
            1'h0:
                casez (\$344 )
                  1'h1:
                      casez (\$350 )
                        1'h1:
                            \fsm_state$next  = 2'h1;
                      endcase
                endcase
            1'h?:
                casez (\$358 )
                  1'h1:
                      casez (\$364 )
                        1'h1:
                            \fsm_state$next  = 2'h1;
                      endcase
                endcase
          endcase
      2'h1:
          casez (\$368 )
            1'h1:
                casez (\$371 )
                  1'h0:
                      casez (\$373 )
                        1'h1:
                            \fsm_state$next  = 2'h2;
                        default:
                            \fsm_state$next  = 2'h3;
                      endcase
                  1'h?:
                      casez (\$375 )
                        1'h1:
                            \fsm_state$next  = 2'h2;
                        default:
                            \fsm_state$next  = 2'h3;
                      endcase
                endcase
          endcase
      2'h2:
          casez (\ready$4 )
            1'h1:
                casez (\$379 )
                  1'h0:
                      casez (\$383 )
                        1'h1:
                            \fsm_state$next  = 2'h3;
                      endcase
                  1'h?:
                      casez (\$387 )
                        1'h1:
                            \fsm_state$next  = 2'h3;
                      endcase
                endcase
          endcase
      2'h3:
        begin
          casez (ack)
            1'h1:
                casez (\$389 )
                  1'h0:
                      casez (buffer_toggle)
                        1'h0:
                            casez ({ \$415 , \$403  })
                              2'b?1:
                                  \fsm_state$next  = 2'h1;
                              2'b1?:
                                  \fsm_state$next  = 2'h1;
                              default:
                                  \fsm_state$next  = 2'h0;
                            endcase
                        1'h?:
                            casez ({ \$433 , \$421  })
                              2'b?1:
                                  \fsm_state$next  = 2'h1;
                              2'b1?:
                                  \fsm_state$next  = 2'h1;
                              default:
                                  \fsm_state$next  = 2'h0;
                            endcase
                      endcase
                  1'h?:
                      casez (buffer_toggle)
                        1'h0:
                            casez ({ \$459 , \$447  })
                              2'b?1:
                                  \fsm_state$next  = 2'h1;
                              2'b1?:
                                  \fsm_state$next  = 2'h1;
                              default:
                                  \fsm_state$next  = 2'h0;
                            endcase
                        1'h?:
                            casez ({ \$477 , \$465  })
                              2'b?1:
                                  \fsm_state$next  = 2'h1;
                              2'b1?:
                                  \fsm_state$next  = 2'h1;
                              default:
                                  \fsm_state$next  = 2'h0;
                            endcase
                      endcase
                endcase
          endcase
          casez (new_token)
            1'h1:
                \fsm_state$next  = 2'h1;
          endcase
        end
    endcase
    casez (usb_rst)
      1'h1:
          \fsm_state$next  = 2'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$31 ) begin end
    \buffer_toggle$next  = buffer_toggle;
    casez (fsm_state)
      2'h0:
          casez (buffer_toggle)
            1'h0:
                casez (\$485 )
                  1'h1:
                      casez (\$491 )
                        1'h1:
                            \buffer_toggle$next  = \$493 ;
                      endcase
                endcase
            1'h?:
                casez (\$501 )
                  1'h1:
                      casez (\$507 )
                        1'h1:
                            \buffer_toggle$next  = \$509 ;
                      endcase
                endcase
          endcase
      2'h1:
          ;
      2'h2:
          ;
      2'h3:
          casez (ack)
            1'h1:
                casez (\$511 )
                  1'h0:
                      casez (buffer_toggle)
                        1'h0:
                            casez ({ \$537 , \$525  })
                              2'b?1:
                                  ;
                              2'b1?:
                                  \buffer_toggle$next  = 1'h0;
                            endcase
                        1'h?:
                            casez ({ \$555 , \$543  })
                              2'b?1:
                                  ;
                              2'b1?:
                                  \buffer_toggle$next  = 1'h0;
                            endcase
                      endcase
                  1'h?:
                      casez (buffer_toggle)
                        1'h0:
                            casez ({ \$581 , \$569  })
                              2'b?1:
                                  ;
                              2'b1?:
                                  \buffer_toggle$next  = 1'h1;
                            endcase
                        1'h?:
                            casez ({ \$599 , \$587  })
                              2'b?1:
                                  ;
                              2'b1?:
                                  \buffer_toggle$next  = 1'h1;
                            endcase
                      endcase
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \buffer_toggle$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$31 ) begin end
    \send_position$next  = send_position;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          \send_position$next  = 10'h000;
      2'h2:
          casez (\ready$4 )
            1'h1:
                \send_position$next  = \$602 [9:0];
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \send_position$next  = 10'h000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$31 ) begin end
    \first$next  = first;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          casez (\$606 )
            1'h1:
                casez (\$609 )
                  1'h0:
                      casez (\$611 )
                        1'h1:
                            \first$next  = 1'h1;
                      endcase
                  1'h?:
                      casez (\$613 )
                        1'h1:
                            \first$next  = 1'h1;
                      endcase
                endcase
          endcase
      2'h2:
          casez (\ready$4 )
            1'h1:
                \first$next  = 1'h0;
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \first$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$31 ) begin end
    casez (buffer_toggle)
      1'h0:
          transmit_buffer_0_w_addr = \$signal [8:0];
      1'h?:
          transmit_buffer_0_w_addr = \$signal$27 [8:0];
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$31 ) begin end
    \valid$1  = 1'h0;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          casez (\$617 )
            1'h1:
                casez (\$620 )
                  1'h0:
                      casez (\$622 )
                        1'h1:
                            ;
                        default:
                            \valid$1  = 1'h1;
                      endcase
                  1'h?:
                      casez (\$624 )
                        1'h1:
                            ;
                        default:
                            \valid$1  = 1'h1;
                      endcase
                endcase
          endcase
      2'h2:
          \valid$1  = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$31 ) begin end
    \last$2  = 1'h0;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          casez (\$628 )
            1'h1:
                casez (\$631 )
                  1'h0:
                      casez (\$633 )
                        1'h1:
                            ;
                        default:
                            \last$2  = 1'h1;
                      endcase
                  1'h?:
                      casez (\$635 )
                        1'h1:
                            ;
                        default:
                            \last$2  = 1'h1;
                      endcase
                endcase
          endcase
      2'h2:
          casez (\$639 )
            1'h0:
                \last$2  = \$643 ;
            1'h?:
                \last$2  = \$647 ;
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$31 ) begin end
    casez (buffer_toggle)
      1'h0:
          transmit_buffer_1_w_addr = \$signal [8:0];
      1'h?:
          transmit_buffer_1_w_addr = \$signal$27 [8:0];
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$31 ) begin end
    transmit_buffer_0_r_addr = 9'h000;
    transmit_buffer_1_r_addr = 9'h000;
    casez (\$156 )
      1'h0:
          transmit_buffer_0_r_addr = send_position[8:0];
      1'h?:
          transmit_buffer_1_r_addr = send_position[8:0];
    endcase
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          ;
      2'h2:
          casez (\ready$4 )
            1'h1:
                casez (\$161 )
                  1'h0:
                      transmit_buffer_0_r_addr = \$164 [8:0];
                  1'h?:
                      transmit_buffer_1_r_addr = \$167 [8:0];
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$31 ) begin end
    casez (\$169 )
      1'h0:
          \payload$3  = transmit_buffer_0_r_data;
      1'h?:
          \payload$3  = transmit_buffer_1_r_data;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$31 ) begin end
    casez (buffer_toggle)
      1'h0:
          ready = \$175 ;
      1'h?:
          ready = \$181 ;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$31 ) begin end
    transmit_buffer_0_w_en = 1'h0;
    transmit_buffer_1_w_en = 1'h0;
    casez (buffer_toggle)
      1'h0:
          transmit_buffer_0_w_en = \$185 ;
      1'h?:
          transmit_buffer_1_w_en = \$187 ;
    endcase
  end
  assign \$151  = \$signal ;
  assign \$152  = \$signal$27 ;
  assign \$154  = \$signal ;
  assign \$155  = \$signal$27 ;
  assign \$158  = \$159 ;
  assign \$163  = \$164 ;
  assign \$166  = \$167 ;
  assign \$189  = \$190 ;
  assign \$192  = \$193 ;
  assign \$601  = \$602 ;
  assign reset_sequence = 1'h0;
  assign start_with_data1 = 1'h0;
  assign transmit_buffer_1_w_data = payload;
  assign transmit_buffer_0_w_data = payload;
  assign \$8  = 1'h1;
  assign \$7  = 2'h1;
  assign \$215  = 1'h1;
  assign \$231  = 1'h0;
  assign \$493  = 1'h1;
  assign \$509  = 1'h0;
endmodule
module \tx_manager$5 (usb_clk, generate_zlps, active, valid, last, payload, ready, \valid$1 , first, \last$2 , \payload$3 , \ready$4 , data_pid, new_token, ready_for_response, is_in, nak, ack, usb_rst);
  reg \$auto$verilog_backend.cc:2083:dump_module$32  = 0;
  wire \$100 ;
  wire \$102 ;
  wire \$104 ;
  wire \$106 ;
  wire \$108 ;
  wire [10:0] \$11 ;
  wire \$110 ;
  wire \$112 ;
  wire [10:0] \$114 ;
  wire \$116 ;
  wire \$118 ;
  wire \$120 ;
  wire \$122 ;
  wire \$124 ;
  wire \$126 ;
  wire \$128 ;
  wire \$13 ;
  wire \$130 ;
  wire \$132 ;
  wire \$134 ;
  wire [10:0] \$136 ;
  wire \$138 ;
  wire \$140 ;
  wire \$142 ;
  wire \$144 ;
  wire \$146 ;
  wire \$148 ;
  wire \$15 ;
  wire [9:0] \$150 ;
  wire [9:0] \$151 ;
  wire [9:0] \$152 ;
  wire [9:0] \$153 ;
  wire [9:0] \$154 ;
  wire [9:0] \$155 ;
  wire \$156 ;
  wire [10:0] \$158 ;
  wire [10:0] \$159 ;
  wire \$161 ;
  wire [10:0] \$163 ;
  wire [10:0] \$164 ;
  wire [10:0] \$166 ;
  wire [10:0] \$167 ;
  wire \$169 ;
  wire \$17 ;
  wire \$171 ;
  wire \$173 ;
  wire \$175 ;
  wire \$177 ;
  wire \$179 ;
  wire \$181 ;
  wire \$183 ;
  wire \$185 ;
  wire \$187 ;
  wire [10:0] \$189 ;
  wire [10:0] \$19 ;
  wire [10:0] \$190 ;
  wire [10:0] \$192 ;
  wire [10:0] \$193 ;
  wire \$195 ;
  wire \$197 ;
  wire \$199 ;
  wire [10:0] \$201 ;
  wire \$203 ;
  wire \$205 ;
  wire \$207 ;
  wire [10:0] \$209 ;
  wire \$21 ;
  wire \$211 ;
  wire \$213 ;
  wire \$215 ;
  wire [10:0] \$217 ;
  wire \$219 ;
  wire \$221 ;
  wire \$223 ;
  wire [10:0] \$225 ;
  wire \$227 ;
  wire \$229 ;
  wire \$23 ;
  wire \$231 ;
  wire \$233 ;
  wire \$235 ;
  wire \$237 ;
  wire \$238 ;
  wire \$240 ;
  wire \$242 ;
  wire \$244 ;
  wire \$246 ;
  wire \$248 ;
  wire \$25 ;
  wire \$250 ;
  wire \$252 ;
  wire \$254 ;
  wire \$256 ;
  wire \$258 ;
  wire \$260 ;
  wire [10:0] \$262 ;
  wire \$264 ;
  wire \$266 ;
  wire \$268 ;
  wire \$270 ;
  wire \$272 ;
  wire \$274 ;
  wire \$276 ;
  wire \$278 ;
  wire [10:0] \$28 ;
  wire [10:0] \$280 ;
  wire \$282 ;
  wire \$284 ;
  wire \$286 ;
  wire \$288 ;
  wire \$290 ;
  wire \$292 ;
  wire \$294 ;
  wire \$296 ;
  wire \$298 ;
  wire \$30 ;
  wire \$300 ;
  wire \$302 ;
  wire \$304 ;
  wire [10:0] \$306 ;
  wire \$308 ;
  wire \$310 ;
  wire \$312 ;
  wire \$314 ;
  wire \$316 ;
  wire \$318 ;
  wire \$32 ;
  wire \$320 ;
  wire \$322 ;
  wire [10:0] \$324 ;
  wire \$326 ;
  wire \$328 ;
  wire \$330 ;
  wire \$332 ;
  wire \$334 ;
  wire \$336 ;
  wire [10:0] \$338 ;
  wire \$34 ;
  wire \$340 ;
  wire \$342 ;
  wire \$344 ;
  wire [10:0] \$346 ;
  wire \$348 ;
  wire \$350 ;
  wire [10:0] \$352 ;
  wire \$354 ;
  wire \$356 ;
  wire \$358 ;
  wire [10:0] \$36 ;
  wire [10:0] \$360 ;
  wire \$362 ;
  wire \$364 ;
  wire \$366 ;
  wire \$368 ;
  wire \$370 ;
  wire \$371 ;
  wire \$373 ;
  wire \$375 ;
  wire [10:0] \$377 ;
  wire \$379 ;
  wire \$38 ;
  wire [10:0] \$381 ;
  wire \$383 ;
  wire [10:0] \$385 ;
  wire \$387 ;
  wire \$389 ;
  wire \$391 ;
  wire \$393 ;
  wire \$395 ;
  wire \$397 ;
  wire \$399 ;
  wire \$40 ;
  wire \$401 ;
  wire \$403 ;
  wire \$405 ;
  wire [10:0] \$407 ;
  wire \$409 ;
  wire \$411 ;
  wire \$413 ;
  wire \$415 ;
  wire \$417 ;
  wire \$419 ;
  wire \$42 ;
  wire \$421 ;
  wire \$423 ;
  wire [10:0] \$425 ;
  wire \$427 ;
  wire \$429 ;
  wire \$431 ;
  wire \$433 ;
  wire \$435 ;
  wire \$437 ;
  wire \$439 ;
  wire \$44 ;
  wire \$441 ;
  wire \$443 ;
  wire \$445 ;
  wire \$447 ;
  wire \$449 ;
  wire [10:0] \$451 ;
  wire \$453 ;
  wire \$455 ;
  wire \$457 ;
  wire \$459 ;
  wire \$46 ;
  wire \$461 ;
  wire \$463 ;
  wire \$465 ;
  wire \$467 ;
  wire [10:0] \$469 ;
  wire \$471 ;
  wire \$473 ;
  wire \$475 ;
  wire \$477 ;
  wire [10:0] \$479 ;
  wire \$48 ;
  wire \$481 ;
  wire \$483 ;
  wire \$485 ;
  wire [10:0] \$487 ;
  wire \$489 ;
  wire \$491 ;
  wire \$493 ;
  wire [10:0] \$495 ;
  wire \$497 ;
  wire \$499 ;
  wire \$50 ;
  wire \$501 ;
  wire [10:0] \$503 ;
  wire \$505 ;
  wire \$507 ;
  wire \$509 ;
  wire \$511 ;
  wire \$513 ;
  wire \$515 ;
  wire \$517 ;
  wire \$519 ;
  wire \$52 ;
  wire \$521 ;
  wire \$523 ;
  wire \$525 ;
  wire \$527 ;
  wire [10:0] \$529 ;
  wire \$531 ;
  wire \$533 ;
  wire \$535 ;
  wire \$537 ;
  wire \$539 ;
  wire \$54 ;
  wire \$541 ;
  wire \$543 ;
  wire \$545 ;
  wire [10:0] \$547 ;
  wire \$549 ;
  wire \$551 ;
  wire \$553 ;
  wire \$555 ;
  wire \$557 ;
  wire \$559 ;
  wire \$56 ;
  wire \$561 ;
  wire \$563 ;
  wire \$565 ;
  wire \$567 ;
  wire \$569 ;
  wire \$571 ;
  wire [10:0] \$573 ;
  wire \$575 ;
  wire \$577 ;
  wire \$579 ;
  wire \$58 ;
  wire \$581 ;
  wire \$583 ;
  wire \$585 ;
  wire \$587 ;
  wire \$589 ;
  wire [10:0] \$591 ;
  wire \$593 ;
  wire \$595 ;
  wire \$597 ;
  wire \$599 ;
  wire \$60 ;
  wire [10:0] \$601 ;
  wire [10:0] \$602 ;
  wire \$604 ;
  wire \$606 ;
  wire \$608 ;
  wire \$609 ;
  wire \$611 ;
  wire \$613 ;
  wire \$615 ;
  wire \$617 ;
  wire \$619 ;
  wire [10:0] \$62 ;
  wire \$620 ;
  wire \$622 ;
  wire \$624 ;
  wire \$626 ;
  wire \$628 ;
  wire \$630 ;
  wire \$631 ;
  wire \$633 ;
  wire \$635 ;
  wire [10:0] \$637 ;
  wire \$639 ;
  wire \$64 ;
  wire [10:0] \$641 ;
  wire \$643 ;
  wire [10:0] \$645 ;
  wire \$647 ;
  wire \$66 ;
  wire \$68 ;
  wire [1:0] \$7 ;
  wire \$70 ;
  wire \$72 ;
  wire \$74 ;
  wire \$76 ;
  wire \$78 ;
  wire \$8 ;
  wire \$80 ;
  wire \$82 ;
  wire [10:0] \$84 ;
  wire \$86 ;
  wire \$88 ;
  wire \$90 ;
  wire \$92 ;
  wire \$94 ;
  wire \$96 ;
  wire \$98 ;
  reg [9:0] \$signal  = 10'h000;
  reg [9:0] \$signal$27  = 10'h000;
  reg [9:0] \$signal$27$next ;
  reg [9:0] \$signal$next ;
  input ack;
  wire ack;
  input active;
  wire active;
  reg buffer_toggle = 1'h0;
  reg \buffer_toggle$next ;
  output [1:0] data_pid;
  reg [1:0] data_pid = 2'h1;
  reg [1:0] \data_pid$next ;
  output first;
  reg first = 1'h0;
  reg \first$next ;
  reg [1:0] fsm_state = 2'h0;
  reg [1:0] \fsm_state$next ;
  input generate_zlps;
  wire generate_zlps;
  input is_in;
  wire is_in;
  input last;
  wire last;
  output \last$2 ;
  reg \last$2 ;
  output nak;
  reg nak;
  input new_token;
  wire new_token;
  input [7:0] payload;
  wire [7:0] payload;
  output [7:0] \payload$3 ;
  reg [7:0] \payload$3 ;
  output ready;
  reg ready;
  input \ready$4 ;
  wire \ready$4 ;
  input ready_for_response;
  wire ready_for_response;
  wire reset_sequence;
  reg [9:0] send_position = 10'h000;
  reg [9:0] \send_position$next ;
  wire start_with_data1;
  reg stream_ended_in_buffer0 = 1'h0;
  reg \stream_ended_in_buffer0$next ;
  reg stream_ended_in_buffer1 = 1'h0;
  reg \stream_ended_in_buffer1$next ;
  reg [8:0] transmit_buffer_0_r_addr;
  wire [7:0] transmit_buffer_0_r_data;
  reg [8:0] transmit_buffer_0_w_addr;
  wire [7:0] transmit_buffer_0_w_data;
  reg transmit_buffer_0_w_en;
  reg [8:0] transmit_buffer_1_r_addr;
  wire [7:0] transmit_buffer_1_r_data;
  reg [8:0] transmit_buffer_1_w_addr;
  wire [7:0] transmit_buffer_1_w_data;
  reg transmit_buffer_1_w_en;
  input usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  input valid;
  wire valid;
  output \valid$1 ;
  reg \valid$1 ;
  reg [7:0] transmit_buffer_0 [511:0];
  initial begin
    transmit_buffer_0[0] = 8'h00;
    transmit_buffer_0[1] = 8'h00;
    transmit_buffer_0[2] = 8'h00;
    transmit_buffer_0[3] = 8'h00;
    transmit_buffer_0[4] = 8'h00;
    transmit_buffer_0[5] = 8'h00;
    transmit_buffer_0[6] = 8'h00;
    transmit_buffer_0[7] = 8'h00;
    transmit_buffer_0[8] = 8'h00;
    transmit_buffer_0[9] = 8'h00;
    transmit_buffer_0[10] = 8'h00;
    transmit_buffer_0[11] = 8'h00;
    transmit_buffer_0[12] = 8'h00;
    transmit_buffer_0[13] = 8'h00;
    transmit_buffer_0[14] = 8'h00;
    transmit_buffer_0[15] = 8'h00;
    transmit_buffer_0[16] = 8'h00;
    transmit_buffer_0[17] = 8'h00;
    transmit_buffer_0[18] = 8'h00;
    transmit_buffer_0[19] = 8'h00;
    transmit_buffer_0[20] = 8'h00;
    transmit_buffer_0[21] = 8'h00;
    transmit_buffer_0[22] = 8'h00;
    transmit_buffer_0[23] = 8'h00;
    transmit_buffer_0[24] = 8'h00;
    transmit_buffer_0[25] = 8'h00;
    transmit_buffer_0[26] = 8'h00;
    transmit_buffer_0[27] = 8'h00;
    transmit_buffer_0[28] = 8'h00;
    transmit_buffer_0[29] = 8'h00;
    transmit_buffer_0[30] = 8'h00;
    transmit_buffer_0[31] = 8'h00;
    transmit_buffer_0[32] = 8'h00;
    transmit_buffer_0[33] = 8'h00;
    transmit_buffer_0[34] = 8'h00;
    transmit_buffer_0[35] = 8'h00;
    transmit_buffer_0[36] = 8'h00;
    transmit_buffer_0[37] = 8'h00;
    transmit_buffer_0[38] = 8'h00;
    transmit_buffer_0[39] = 8'h00;
    transmit_buffer_0[40] = 8'h00;
    transmit_buffer_0[41] = 8'h00;
    transmit_buffer_0[42] = 8'h00;
    transmit_buffer_0[43] = 8'h00;
    transmit_buffer_0[44] = 8'h00;
    transmit_buffer_0[45] = 8'h00;
    transmit_buffer_0[46] = 8'h00;
    transmit_buffer_0[47] = 8'h00;
    transmit_buffer_0[48] = 8'h00;
    transmit_buffer_0[49] = 8'h00;
    transmit_buffer_0[50] = 8'h00;
    transmit_buffer_0[51] = 8'h00;
    transmit_buffer_0[52] = 8'h00;
    transmit_buffer_0[53] = 8'h00;
    transmit_buffer_0[54] = 8'h00;
    transmit_buffer_0[55] = 8'h00;
    transmit_buffer_0[56] = 8'h00;
    transmit_buffer_0[57] = 8'h00;
    transmit_buffer_0[58] = 8'h00;
    transmit_buffer_0[59] = 8'h00;
    transmit_buffer_0[60] = 8'h00;
    transmit_buffer_0[61] = 8'h00;
    transmit_buffer_0[62] = 8'h00;
    transmit_buffer_0[63] = 8'h00;
    transmit_buffer_0[64] = 8'h00;
    transmit_buffer_0[65] = 8'h00;
    transmit_buffer_0[66] = 8'h00;
    transmit_buffer_0[67] = 8'h00;
    transmit_buffer_0[68] = 8'h00;
    transmit_buffer_0[69] = 8'h00;
    transmit_buffer_0[70] = 8'h00;
    transmit_buffer_0[71] = 8'h00;
    transmit_buffer_0[72] = 8'h00;
    transmit_buffer_0[73] = 8'h00;
    transmit_buffer_0[74] = 8'h00;
    transmit_buffer_0[75] = 8'h00;
    transmit_buffer_0[76] = 8'h00;
    transmit_buffer_0[77] = 8'h00;
    transmit_buffer_0[78] = 8'h00;
    transmit_buffer_0[79] = 8'h00;
    transmit_buffer_0[80] = 8'h00;
    transmit_buffer_0[81] = 8'h00;
    transmit_buffer_0[82] = 8'h00;
    transmit_buffer_0[83] = 8'h00;
    transmit_buffer_0[84] = 8'h00;
    transmit_buffer_0[85] = 8'h00;
    transmit_buffer_0[86] = 8'h00;
    transmit_buffer_0[87] = 8'h00;
    transmit_buffer_0[88] = 8'h00;
    transmit_buffer_0[89] = 8'h00;
    transmit_buffer_0[90] = 8'h00;
    transmit_buffer_0[91] = 8'h00;
    transmit_buffer_0[92] = 8'h00;
    transmit_buffer_0[93] = 8'h00;
    transmit_buffer_0[94] = 8'h00;
    transmit_buffer_0[95] = 8'h00;
    transmit_buffer_0[96] = 8'h00;
    transmit_buffer_0[97] = 8'h00;
    transmit_buffer_0[98] = 8'h00;
    transmit_buffer_0[99] = 8'h00;
    transmit_buffer_0[100] = 8'h00;
    transmit_buffer_0[101] = 8'h00;
    transmit_buffer_0[102] = 8'h00;
    transmit_buffer_0[103] = 8'h00;
    transmit_buffer_0[104] = 8'h00;
    transmit_buffer_0[105] = 8'h00;
    transmit_buffer_0[106] = 8'h00;
    transmit_buffer_0[107] = 8'h00;
    transmit_buffer_0[108] = 8'h00;
    transmit_buffer_0[109] = 8'h00;
    transmit_buffer_0[110] = 8'h00;
    transmit_buffer_0[111] = 8'h00;
    transmit_buffer_0[112] = 8'h00;
    transmit_buffer_0[113] = 8'h00;
    transmit_buffer_0[114] = 8'h00;
    transmit_buffer_0[115] = 8'h00;
    transmit_buffer_0[116] = 8'h00;
    transmit_buffer_0[117] = 8'h00;
    transmit_buffer_0[118] = 8'h00;
    transmit_buffer_0[119] = 8'h00;
    transmit_buffer_0[120] = 8'h00;
    transmit_buffer_0[121] = 8'h00;
    transmit_buffer_0[122] = 8'h00;
    transmit_buffer_0[123] = 8'h00;
    transmit_buffer_0[124] = 8'h00;
    transmit_buffer_0[125] = 8'h00;
    transmit_buffer_0[126] = 8'h00;
    transmit_buffer_0[127] = 8'h00;
    transmit_buffer_0[128] = 8'h00;
    transmit_buffer_0[129] = 8'h00;
    transmit_buffer_0[130] = 8'h00;
    transmit_buffer_0[131] = 8'h00;
    transmit_buffer_0[132] = 8'h00;
    transmit_buffer_0[133] = 8'h00;
    transmit_buffer_0[134] = 8'h00;
    transmit_buffer_0[135] = 8'h00;
    transmit_buffer_0[136] = 8'h00;
    transmit_buffer_0[137] = 8'h00;
    transmit_buffer_0[138] = 8'h00;
    transmit_buffer_0[139] = 8'h00;
    transmit_buffer_0[140] = 8'h00;
    transmit_buffer_0[141] = 8'h00;
    transmit_buffer_0[142] = 8'h00;
    transmit_buffer_0[143] = 8'h00;
    transmit_buffer_0[144] = 8'h00;
    transmit_buffer_0[145] = 8'h00;
    transmit_buffer_0[146] = 8'h00;
    transmit_buffer_0[147] = 8'h00;
    transmit_buffer_0[148] = 8'h00;
    transmit_buffer_0[149] = 8'h00;
    transmit_buffer_0[150] = 8'h00;
    transmit_buffer_0[151] = 8'h00;
    transmit_buffer_0[152] = 8'h00;
    transmit_buffer_0[153] = 8'h00;
    transmit_buffer_0[154] = 8'h00;
    transmit_buffer_0[155] = 8'h00;
    transmit_buffer_0[156] = 8'h00;
    transmit_buffer_0[157] = 8'h00;
    transmit_buffer_0[158] = 8'h00;
    transmit_buffer_0[159] = 8'h00;
    transmit_buffer_0[160] = 8'h00;
    transmit_buffer_0[161] = 8'h00;
    transmit_buffer_0[162] = 8'h00;
    transmit_buffer_0[163] = 8'h00;
    transmit_buffer_0[164] = 8'h00;
    transmit_buffer_0[165] = 8'h00;
    transmit_buffer_0[166] = 8'h00;
    transmit_buffer_0[167] = 8'h00;
    transmit_buffer_0[168] = 8'h00;
    transmit_buffer_0[169] = 8'h00;
    transmit_buffer_0[170] = 8'h00;
    transmit_buffer_0[171] = 8'h00;
    transmit_buffer_0[172] = 8'h00;
    transmit_buffer_0[173] = 8'h00;
    transmit_buffer_0[174] = 8'h00;
    transmit_buffer_0[175] = 8'h00;
    transmit_buffer_0[176] = 8'h00;
    transmit_buffer_0[177] = 8'h00;
    transmit_buffer_0[178] = 8'h00;
    transmit_buffer_0[179] = 8'h00;
    transmit_buffer_0[180] = 8'h00;
    transmit_buffer_0[181] = 8'h00;
    transmit_buffer_0[182] = 8'h00;
    transmit_buffer_0[183] = 8'h00;
    transmit_buffer_0[184] = 8'h00;
    transmit_buffer_0[185] = 8'h00;
    transmit_buffer_0[186] = 8'h00;
    transmit_buffer_0[187] = 8'h00;
    transmit_buffer_0[188] = 8'h00;
    transmit_buffer_0[189] = 8'h00;
    transmit_buffer_0[190] = 8'h00;
    transmit_buffer_0[191] = 8'h00;
    transmit_buffer_0[192] = 8'h00;
    transmit_buffer_0[193] = 8'h00;
    transmit_buffer_0[194] = 8'h00;
    transmit_buffer_0[195] = 8'h00;
    transmit_buffer_0[196] = 8'h00;
    transmit_buffer_0[197] = 8'h00;
    transmit_buffer_0[198] = 8'h00;
    transmit_buffer_0[199] = 8'h00;
    transmit_buffer_0[200] = 8'h00;
    transmit_buffer_0[201] = 8'h00;
    transmit_buffer_0[202] = 8'h00;
    transmit_buffer_0[203] = 8'h00;
    transmit_buffer_0[204] = 8'h00;
    transmit_buffer_0[205] = 8'h00;
    transmit_buffer_0[206] = 8'h00;
    transmit_buffer_0[207] = 8'h00;
    transmit_buffer_0[208] = 8'h00;
    transmit_buffer_0[209] = 8'h00;
    transmit_buffer_0[210] = 8'h00;
    transmit_buffer_0[211] = 8'h00;
    transmit_buffer_0[212] = 8'h00;
    transmit_buffer_0[213] = 8'h00;
    transmit_buffer_0[214] = 8'h00;
    transmit_buffer_0[215] = 8'h00;
    transmit_buffer_0[216] = 8'h00;
    transmit_buffer_0[217] = 8'h00;
    transmit_buffer_0[218] = 8'h00;
    transmit_buffer_0[219] = 8'h00;
    transmit_buffer_0[220] = 8'h00;
    transmit_buffer_0[221] = 8'h00;
    transmit_buffer_0[222] = 8'h00;
    transmit_buffer_0[223] = 8'h00;
    transmit_buffer_0[224] = 8'h00;
    transmit_buffer_0[225] = 8'h00;
    transmit_buffer_0[226] = 8'h00;
    transmit_buffer_0[227] = 8'h00;
    transmit_buffer_0[228] = 8'h00;
    transmit_buffer_0[229] = 8'h00;
    transmit_buffer_0[230] = 8'h00;
    transmit_buffer_0[231] = 8'h00;
    transmit_buffer_0[232] = 8'h00;
    transmit_buffer_0[233] = 8'h00;
    transmit_buffer_0[234] = 8'h00;
    transmit_buffer_0[235] = 8'h00;
    transmit_buffer_0[236] = 8'h00;
    transmit_buffer_0[237] = 8'h00;
    transmit_buffer_0[238] = 8'h00;
    transmit_buffer_0[239] = 8'h00;
    transmit_buffer_0[240] = 8'h00;
    transmit_buffer_0[241] = 8'h00;
    transmit_buffer_0[242] = 8'h00;
    transmit_buffer_0[243] = 8'h00;
    transmit_buffer_0[244] = 8'h00;
    transmit_buffer_0[245] = 8'h00;
    transmit_buffer_0[246] = 8'h00;
    transmit_buffer_0[247] = 8'h00;
    transmit_buffer_0[248] = 8'h00;
    transmit_buffer_0[249] = 8'h00;
    transmit_buffer_0[250] = 8'h00;
    transmit_buffer_0[251] = 8'h00;
    transmit_buffer_0[252] = 8'h00;
    transmit_buffer_0[253] = 8'h00;
    transmit_buffer_0[254] = 8'h00;
    transmit_buffer_0[255] = 8'h00;
    transmit_buffer_0[256] = 8'h00;
    transmit_buffer_0[257] = 8'h00;
    transmit_buffer_0[258] = 8'h00;
    transmit_buffer_0[259] = 8'h00;
    transmit_buffer_0[260] = 8'h00;
    transmit_buffer_0[261] = 8'h00;
    transmit_buffer_0[262] = 8'h00;
    transmit_buffer_0[263] = 8'h00;
    transmit_buffer_0[264] = 8'h00;
    transmit_buffer_0[265] = 8'h00;
    transmit_buffer_0[266] = 8'h00;
    transmit_buffer_0[267] = 8'h00;
    transmit_buffer_0[268] = 8'h00;
    transmit_buffer_0[269] = 8'h00;
    transmit_buffer_0[270] = 8'h00;
    transmit_buffer_0[271] = 8'h00;
    transmit_buffer_0[272] = 8'h00;
    transmit_buffer_0[273] = 8'h00;
    transmit_buffer_0[274] = 8'h00;
    transmit_buffer_0[275] = 8'h00;
    transmit_buffer_0[276] = 8'h00;
    transmit_buffer_0[277] = 8'h00;
    transmit_buffer_0[278] = 8'h00;
    transmit_buffer_0[279] = 8'h00;
    transmit_buffer_0[280] = 8'h00;
    transmit_buffer_0[281] = 8'h00;
    transmit_buffer_0[282] = 8'h00;
    transmit_buffer_0[283] = 8'h00;
    transmit_buffer_0[284] = 8'h00;
    transmit_buffer_0[285] = 8'h00;
    transmit_buffer_0[286] = 8'h00;
    transmit_buffer_0[287] = 8'h00;
    transmit_buffer_0[288] = 8'h00;
    transmit_buffer_0[289] = 8'h00;
    transmit_buffer_0[290] = 8'h00;
    transmit_buffer_0[291] = 8'h00;
    transmit_buffer_0[292] = 8'h00;
    transmit_buffer_0[293] = 8'h00;
    transmit_buffer_0[294] = 8'h00;
    transmit_buffer_0[295] = 8'h00;
    transmit_buffer_0[296] = 8'h00;
    transmit_buffer_0[297] = 8'h00;
    transmit_buffer_0[298] = 8'h00;
    transmit_buffer_0[299] = 8'h00;
    transmit_buffer_0[300] = 8'h00;
    transmit_buffer_0[301] = 8'h00;
    transmit_buffer_0[302] = 8'h00;
    transmit_buffer_0[303] = 8'h00;
    transmit_buffer_0[304] = 8'h00;
    transmit_buffer_0[305] = 8'h00;
    transmit_buffer_0[306] = 8'h00;
    transmit_buffer_0[307] = 8'h00;
    transmit_buffer_0[308] = 8'h00;
    transmit_buffer_0[309] = 8'h00;
    transmit_buffer_0[310] = 8'h00;
    transmit_buffer_0[311] = 8'h00;
    transmit_buffer_0[312] = 8'h00;
    transmit_buffer_0[313] = 8'h00;
    transmit_buffer_0[314] = 8'h00;
    transmit_buffer_0[315] = 8'h00;
    transmit_buffer_0[316] = 8'h00;
    transmit_buffer_0[317] = 8'h00;
    transmit_buffer_0[318] = 8'h00;
    transmit_buffer_0[319] = 8'h00;
    transmit_buffer_0[320] = 8'h00;
    transmit_buffer_0[321] = 8'h00;
    transmit_buffer_0[322] = 8'h00;
    transmit_buffer_0[323] = 8'h00;
    transmit_buffer_0[324] = 8'h00;
    transmit_buffer_0[325] = 8'h00;
    transmit_buffer_0[326] = 8'h00;
    transmit_buffer_0[327] = 8'h00;
    transmit_buffer_0[328] = 8'h00;
    transmit_buffer_0[329] = 8'h00;
    transmit_buffer_0[330] = 8'h00;
    transmit_buffer_0[331] = 8'h00;
    transmit_buffer_0[332] = 8'h00;
    transmit_buffer_0[333] = 8'h00;
    transmit_buffer_0[334] = 8'h00;
    transmit_buffer_0[335] = 8'h00;
    transmit_buffer_0[336] = 8'h00;
    transmit_buffer_0[337] = 8'h00;
    transmit_buffer_0[338] = 8'h00;
    transmit_buffer_0[339] = 8'h00;
    transmit_buffer_0[340] = 8'h00;
    transmit_buffer_0[341] = 8'h00;
    transmit_buffer_0[342] = 8'h00;
    transmit_buffer_0[343] = 8'h00;
    transmit_buffer_0[344] = 8'h00;
    transmit_buffer_0[345] = 8'h00;
    transmit_buffer_0[346] = 8'h00;
    transmit_buffer_0[347] = 8'h00;
    transmit_buffer_0[348] = 8'h00;
    transmit_buffer_0[349] = 8'h00;
    transmit_buffer_0[350] = 8'h00;
    transmit_buffer_0[351] = 8'h00;
    transmit_buffer_0[352] = 8'h00;
    transmit_buffer_0[353] = 8'h00;
    transmit_buffer_0[354] = 8'h00;
    transmit_buffer_0[355] = 8'h00;
    transmit_buffer_0[356] = 8'h00;
    transmit_buffer_0[357] = 8'h00;
    transmit_buffer_0[358] = 8'h00;
    transmit_buffer_0[359] = 8'h00;
    transmit_buffer_0[360] = 8'h00;
    transmit_buffer_0[361] = 8'h00;
    transmit_buffer_0[362] = 8'h00;
    transmit_buffer_0[363] = 8'h00;
    transmit_buffer_0[364] = 8'h00;
    transmit_buffer_0[365] = 8'h00;
    transmit_buffer_0[366] = 8'h00;
    transmit_buffer_0[367] = 8'h00;
    transmit_buffer_0[368] = 8'h00;
    transmit_buffer_0[369] = 8'h00;
    transmit_buffer_0[370] = 8'h00;
    transmit_buffer_0[371] = 8'h00;
    transmit_buffer_0[372] = 8'h00;
    transmit_buffer_0[373] = 8'h00;
    transmit_buffer_0[374] = 8'h00;
    transmit_buffer_0[375] = 8'h00;
    transmit_buffer_0[376] = 8'h00;
    transmit_buffer_0[377] = 8'h00;
    transmit_buffer_0[378] = 8'h00;
    transmit_buffer_0[379] = 8'h00;
    transmit_buffer_0[380] = 8'h00;
    transmit_buffer_0[381] = 8'h00;
    transmit_buffer_0[382] = 8'h00;
    transmit_buffer_0[383] = 8'h00;
    transmit_buffer_0[384] = 8'h00;
    transmit_buffer_0[385] = 8'h00;
    transmit_buffer_0[386] = 8'h00;
    transmit_buffer_0[387] = 8'h00;
    transmit_buffer_0[388] = 8'h00;
    transmit_buffer_0[389] = 8'h00;
    transmit_buffer_0[390] = 8'h00;
    transmit_buffer_0[391] = 8'h00;
    transmit_buffer_0[392] = 8'h00;
    transmit_buffer_0[393] = 8'h00;
    transmit_buffer_0[394] = 8'h00;
    transmit_buffer_0[395] = 8'h00;
    transmit_buffer_0[396] = 8'h00;
    transmit_buffer_0[397] = 8'h00;
    transmit_buffer_0[398] = 8'h00;
    transmit_buffer_0[399] = 8'h00;
    transmit_buffer_0[400] = 8'h00;
    transmit_buffer_0[401] = 8'h00;
    transmit_buffer_0[402] = 8'h00;
    transmit_buffer_0[403] = 8'h00;
    transmit_buffer_0[404] = 8'h00;
    transmit_buffer_0[405] = 8'h00;
    transmit_buffer_0[406] = 8'h00;
    transmit_buffer_0[407] = 8'h00;
    transmit_buffer_0[408] = 8'h00;
    transmit_buffer_0[409] = 8'h00;
    transmit_buffer_0[410] = 8'h00;
    transmit_buffer_0[411] = 8'h00;
    transmit_buffer_0[412] = 8'h00;
    transmit_buffer_0[413] = 8'h00;
    transmit_buffer_0[414] = 8'h00;
    transmit_buffer_0[415] = 8'h00;
    transmit_buffer_0[416] = 8'h00;
    transmit_buffer_0[417] = 8'h00;
    transmit_buffer_0[418] = 8'h00;
    transmit_buffer_0[419] = 8'h00;
    transmit_buffer_0[420] = 8'h00;
    transmit_buffer_0[421] = 8'h00;
    transmit_buffer_0[422] = 8'h00;
    transmit_buffer_0[423] = 8'h00;
    transmit_buffer_0[424] = 8'h00;
    transmit_buffer_0[425] = 8'h00;
    transmit_buffer_0[426] = 8'h00;
    transmit_buffer_0[427] = 8'h00;
    transmit_buffer_0[428] = 8'h00;
    transmit_buffer_0[429] = 8'h00;
    transmit_buffer_0[430] = 8'h00;
    transmit_buffer_0[431] = 8'h00;
    transmit_buffer_0[432] = 8'h00;
    transmit_buffer_0[433] = 8'h00;
    transmit_buffer_0[434] = 8'h00;
    transmit_buffer_0[435] = 8'h00;
    transmit_buffer_0[436] = 8'h00;
    transmit_buffer_0[437] = 8'h00;
    transmit_buffer_0[438] = 8'h00;
    transmit_buffer_0[439] = 8'h00;
    transmit_buffer_0[440] = 8'h00;
    transmit_buffer_0[441] = 8'h00;
    transmit_buffer_0[442] = 8'h00;
    transmit_buffer_0[443] = 8'h00;
    transmit_buffer_0[444] = 8'h00;
    transmit_buffer_0[445] = 8'h00;
    transmit_buffer_0[446] = 8'h00;
    transmit_buffer_0[447] = 8'h00;
    transmit_buffer_0[448] = 8'h00;
    transmit_buffer_0[449] = 8'h00;
    transmit_buffer_0[450] = 8'h00;
    transmit_buffer_0[451] = 8'h00;
    transmit_buffer_0[452] = 8'h00;
    transmit_buffer_0[453] = 8'h00;
    transmit_buffer_0[454] = 8'h00;
    transmit_buffer_0[455] = 8'h00;
    transmit_buffer_0[456] = 8'h00;
    transmit_buffer_0[457] = 8'h00;
    transmit_buffer_0[458] = 8'h00;
    transmit_buffer_0[459] = 8'h00;
    transmit_buffer_0[460] = 8'h00;
    transmit_buffer_0[461] = 8'h00;
    transmit_buffer_0[462] = 8'h00;
    transmit_buffer_0[463] = 8'h00;
    transmit_buffer_0[464] = 8'h00;
    transmit_buffer_0[465] = 8'h00;
    transmit_buffer_0[466] = 8'h00;
    transmit_buffer_0[467] = 8'h00;
    transmit_buffer_0[468] = 8'h00;
    transmit_buffer_0[469] = 8'h00;
    transmit_buffer_0[470] = 8'h00;
    transmit_buffer_0[471] = 8'h00;
    transmit_buffer_0[472] = 8'h00;
    transmit_buffer_0[473] = 8'h00;
    transmit_buffer_0[474] = 8'h00;
    transmit_buffer_0[475] = 8'h00;
    transmit_buffer_0[476] = 8'h00;
    transmit_buffer_0[477] = 8'h00;
    transmit_buffer_0[478] = 8'h00;
    transmit_buffer_0[479] = 8'h00;
    transmit_buffer_0[480] = 8'h00;
    transmit_buffer_0[481] = 8'h00;
    transmit_buffer_0[482] = 8'h00;
    transmit_buffer_0[483] = 8'h00;
    transmit_buffer_0[484] = 8'h00;
    transmit_buffer_0[485] = 8'h00;
    transmit_buffer_0[486] = 8'h00;
    transmit_buffer_0[487] = 8'h00;
    transmit_buffer_0[488] = 8'h00;
    transmit_buffer_0[489] = 8'h00;
    transmit_buffer_0[490] = 8'h00;
    transmit_buffer_0[491] = 8'h00;
    transmit_buffer_0[492] = 8'h00;
    transmit_buffer_0[493] = 8'h00;
    transmit_buffer_0[494] = 8'h00;
    transmit_buffer_0[495] = 8'h00;
    transmit_buffer_0[496] = 8'h00;
    transmit_buffer_0[497] = 8'h00;
    transmit_buffer_0[498] = 8'h00;
    transmit_buffer_0[499] = 8'h00;
    transmit_buffer_0[500] = 8'h00;
    transmit_buffer_0[501] = 8'h00;
    transmit_buffer_0[502] = 8'h00;
    transmit_buffer_0[503] = 8'h00;
    transmit_buffer_0[504] = 8'h00;
    transmit_buffer_0[505] = 8'h00;
    transmit_buffer_0[506] = 8'h00;
    transmit_buffer_0[507] = 8'h00;
    transmit_buffer_0[508] = 8'h00;
    transmit_buffer_0[509] = 8'h00;
    transmit_buffer_0[510] = 8'h00;
    transmit_buffer_0[511] = 8'h00;
  end
  always @(posedge usb_clk) begin
    if (transmit_buffer_0_w_en)
      transmit_buffer_0[transmit_buffer_0_w_addr] <= transmit_buffer_0_w_data;
  end
  reg [8:0] _0_;
  always @(posedge usb_clk) begin
    _0_ <= transmit_buffer_0_r_addr;
  end
  assign transmit_buffer_0_r_data = transmit_buffer_0[_0_];
  reg [7:0] transmit_buffer_1 [511:0];
  initial begin
    transmit_buffer_1[0] = 8'h00;
    transmit_buffer_1[1] = 8'h00;
    transmit_buffer_1[2] = 8'h00;
    transmit_buffer_1[3] = 8'h00;
    transmit_buffer_1[4] = 8'h00;
    transmit_buffer_1[5] = 8'h00;
    transmit_buffer_1[6] = 8'h00;
    transmit_buffer_1[7] = 8'h00;
    transmit_buffer_1[8] = 8'h00;
    transmit_buffer_1[9] = 8'h00;
    transmit_buffer_1[10] = 8'h00;
    transmit_buffer_1[11] = 8'h00;
    transmit_buffer_1[12] = 8'h00;
    transmit_buffer_1[13] = 8'h00;
    transmit_buffer_1[14] = 8'h00;
    transmit_buffer_1[15] = 8'h00;
    transmit_buffer_1[16] = 8'h00;
    transmit_buffer_1[17] = 8'h00;
    transmit_buffer_1[18] = 8'h00;
    transmit_buffer_1[19] = 8'h00;
    transmit_buffer_1[20] = 8'h00;
    transmit_buffer_1[21] = 8'h00;
    transmit_buffer_1[22] = 8'h00;
    transmit_buffer_1[23] = 8'h00;
    transmit_buffer_1[24] = 8'h00;
    transmit_buffer_1[25] = 8'h00;
    transmit_buffer_1[26] = 8'h00;
    transmit_buffer_1[27] = 8'h00;
    transmit_buffer_1[28] = 8'h00;
    transmit_buffer_1[29] = 8'h00;
    transmit_buffer_1[30] = 8'h00;
    transmit_buffer_1[31] = 8'h00;
    transmit_buffer_1[32] = 8'h00;
    transmit_buffer_1[33] = 8'h00;
    transmit_buffer_1[34] = 8'h00;
    transmit_buffer_1[35] = 8'h00;
    transmit_buffer_1[36] = 8'h00;
    transmit_buffer_1[37] = 8'h00;
    transmit_buffer_1[38] = 8'h00;
    transmit_buffer_1[39] = 8'h00;
    transmit_buffer_1[40] = 8'h00;
    transmit_buffer_1[41] = 8'h00;
    transmit_buffer_1[42] = 8'h00;
    transmit_buffer_1[43] = 8'h00;
    transmit_buffer_1[44] = 8'h00;
    transmit_buffer_1[45] = 8'h00;
    transmit_buffer_1[46] = 8'h00;
    transmit_buffer_1[47] = 8'h00;
    transmit_buffer_1[48] = 8'h00;
    transmit_buffer_1[49] = 8'h00;
    transmit_buffer_1[50] = 8'h00;
    transmit_buffer_1[51] = 8'h00;
    transmit_buffer_1[52] = 8'h00;
    transmit_buffer_1[53] = 8'h00;
    transmit_buffer_1[54] = 8'h00;
    transmit_buffer_1[55] = 8'h00;
    transmit_buffer_1[56] = 8'h00;
    transmit_buffer_1[57] = 8'h00;
    transmit_buffer_1[58] = 8'h00;
    transmit_buffer_1[59] = 8'h00;
    transmit_buffer_1[60] = 8'h00;
    transmit_buffer_1[61] = 8'h00;
    transmit_buffer_1[62] = 8'h00;
    transmit_buffer_1[63] = 8'h00;
    transmit_buffer_1[64] = 8'h00;
    transmit_buffer_1[65] = 8'h00;
    transmit_buffer_1[66] = 8'h00;
    transmit_buffer_1[67] = 8'h00;
    transmit_buffer_1[68] = 8'h00;
    transmit_buffer_1[69] = 8'h00;
    transmit_buffer_1[70] = 8'h00;
    transmit_buffer_1[71] = 8'h00;
    transmit_buffer_1[72] = 8'h00;
    transmit_buffer_1[73] = 8'h00;
    transmit_buffer_1[74] = 8'h00;
    transmit_buffer_1[75] = 8'h00;
    transmit_buffer_1[76] = 8'h00;
    transmit_buffer_1[77] = 8'h00;
    transmit_buffer_1[78] = 8'h00;
    transmit_buffer_1[79] = 8'h00;
    transmit_buffer_1[80] = 8'h00;
    transmit_buffer_1[81] = 8'h00;
    transmit_buffer_1[82] = 8'h00;
    transmit_buffer_1[83] = 8'h00;
    transmit_buffer_1[84] = 8'h00;
    transmit_buffer_1[85] = 8'h00;
    transmit_buffer_1[86] = 8'h00;
    transmit_buffer_1[87] = 8'h00;
    transmit_buffer_1[88] = 8'h00;
    transmit_buffer_1[89] = 8'h00;
    transmit_buffer_1[90] = 8'h00;
    transmit_buffer_1[91] = 8'h00;
    transmit_buffer_1[92] = 8'h00;
    transmit_buffer_1[93] = 8'h00;
    transmit_buffer_1[94] = 8'h00;
    transmit_buffer_1[95] = 8'h00;
    transmit_buffer_1[96] = 8'h00;
    transmit_buffer_1[97] = 8'h00;
    transmit_buffer_1[98] = 8'h00;
    transmit_buffer_1[99] = 8'h00;
    transmit_buffer_1[100] = 8'h00;
    transmit_buffer_1[101] = 8'h00;
    transmit_buffer_1[102] = 8'h00;
    transmit_buffer_1[103] = 8'h00;
    transmit_buffer_1[104] = 8'h00;
    transmit_buffer_1[105] = 8'h00;
    transmit_buffer_1[106] = 8'h00;
    transmit_buffer_1[107] = 8'h00;
    transmit_buffer_1[108] = 8'h00;
    transmit_buffer_1[109] = 8'h00;
    transmit_buffer_1[110] = 8'h00;
    transmit_buffer_1[111] = 8'h00;
    transmit_buffer_1[112] = 8'h00;
    transmit_buffer_1[113] = 8'h00;
    transmit_buffer_1[114] = 8'h00;
    transmit_buffer_1[115] = 8'h00;
    transmit_buffer_1[116] = 8'h00;
    transmit_buffer_1[117] = 8'h00;
    transmit_buffer_1[118] = 8'h00;
    transmit_buffer_1[119] = 8'h00;
    transmit_buffer_1[120] = 8'h00;
    transmit_buffer_1[121] = 8'h00;
    transmit_buffer_1[122] = 8'h00;
    transmit_buffer_1[123] = 8'h00;
    transmit_buffer_1[124] = 8'h00;
    transmit_buffer_1[125] = 8'h00;
    transmit_buffer_1[126] = 8'h00;
    transmit_buffer_1[127] = 8'h00;
    transmit_buffer_1[128] = 8'h00;
    transmit_buffer_1[129] = 8'h00;
    transmit_buffer_1[130] = 8'h00;
    transmit_buffer_1[131] = 8'h00;
    transmit_buffer_1[132] = 8'h00;
    transmit_buffer_1[133] = 8'h00;
    transmit_buffer_1[134] = 8'h00;
    transmit_buffer_1[135] = 8'h00;
    transmit_buffer_1[136] = 8'h00;
    transmit_buffer_1[137] = 8'h00;
    transmit_buffer_1[138] = 8'h00;
    transmit_buffer_1[139] = 8'h00;
    transmit_buffer_1[140] = 8'h00;
    transmit_buffer_1[141] = 8'h00;
    transmit_buffer_1[142] = 8'h00;
    transmit_buffer_1[143] = 8'h00;
    transmit_buffer_1[144] = 8'h00;
    transmit_buffer_1[145] = 8'h00;
    transmit_buffer_1[146] = 8'h00;
    transmit_buffer_1[147] = 8'h00;
    transmit_buffer_1[148] = 8'h00;
    transmit_buffer_1[149] = 8'h00;
    transmit_buffer_1[150] = 8'h00;
    transmit_buffer_1[151] = 8'h00;
    transmit_buffer_1[152] = 8'h00;
    transmit_buffer_1[153] = 8'h00;
    transmit_buffer_1[154] = 8'h00;
    transmit_buffer_1[155] = 8'h00;
    transmit_buffer_1[156] = 8'h00;
    transmit_buffer_1[157] = 8'h00;
    transmit_buffer_1[158] = 8'h00;
    transmit_buffer_1[159] = 8'h00;
    transmit_buffer_1[160] = 8'h00;
    transmit_buffer_1[161] = 8'h00;
    transmit_buffer_1[162] = 8'h00;
    transmit_buffer_1[163] = 8'h00;
    transmit_buffer_1[164] = 8'h00;
    transmit_buffer_1[165] = 8'h00;
    transmit_buffer_1[166] = 8'h00;
    transmit_buffer_1[167] = 8'h00;
    transmit_buffer_1[168] = 8'h00;
    transmit_buffer_1[169] = 8'h00;
    transmit_buffer_1[170] = 8'h00;
    transmit_buffer_1[171] = 8'h00;
    transmit_buffer_1[172] = 8'h00;
    transmit_buffer_1[173] = 8'h00;
    transmit_buffer_1[174] = 8'h00;
    transmit_buffer_1[175] = 8'h00;
    transmit_buffer_1[176] = 8'h00;
    transmit_buffer_1[177] = 8'h00;
    transmit_buffer_1[178] = 8'h00;
    transmit_buffer_1[179] = 8'h00;
    transmit_buffer_1[180] = 8'h00;
    transmit_buffer_1[181] = 8'h00;
    transmit_buffer_1[182] = 8'h00;
    transmit_buffer_1[183] = 8'h00;
    transmit_buffer_1[184] = 8'h00;
    transmit_buffer_1[185] = 8'h00;
    transmit_buffer_1[186] = 8'h00;
    transmit_buffer_1[187] = 8'h00;
    transmit_buffer_1[188] = 8'h00;
    transmit_buffer_1[189] = 8'h00;
    transmit_buffer_1[190] = 8'h00;
    transmit_buffer_1[191] = 8'h00;
    transmit_buffer_1[192] = 8'h00;
    transmit_buffer_1[193] = 8'h00;
    transmit_buffer_1[194] = 8'h00;
    transmit_buffer_1[195] = 8'h00;
    transmit_buffer_1[196] = 8'h00;
    transmit_buffer_1[197] = 8'h00;
    transmit_buffer_1[198] = 8'h00;
    transmit_buffer_1[199] = 8'h00;
    transmit_buffer_1[200] = 8'h00;
    transmit_buffer_1[201] = 8'h00;
    transmit_buffer_1[202] = 8'h00;
    transmit_buffer_1[203] = 8'h00;
    transmit_buffer_1[204] = 8'h00;
    transmit_buffer_1[205] = 8'h00;
    transmit_buffer_1[206] = 8'h00;
    transmit_buffer_1[207] = 8'h00;
    transmit_buffer_1[208] = 8'h00;
    transmit_buffer_1[209] = 8'h00;
    transmit_buffer_1[210] = 8'h00;
    transmit_buffer_1[211] = 8'h00;
    transmit_buffer_1[212] = 8'h00;
    transmit_buffer_1[213] = 8'h00;
    transmit_buffer_1[214] = 8'h00;
    transmit_buffer_1[215] = 8'h00;
    transmit_buffer_1[216] = 8'h00;
    transmit_buffer_1[217] = 8'h00;
    transmit_buffer_1[218] = 8'h00;
    transmit_buffer_1[219] = 8'h00;
    transmit_buffer_1[220] = 8'h00;
    transmit_buffer_1[221] = 8'h00;
    transmit_buffer_1[222] = 8'h00;
    transmit_buffer_1[223] = 8'h00;
    transmit_buffer_1[224] = 8'h00;
    transmit_buffer_1[225] = 8'h00;
    transmit_buffer_1[226] = 8'h00;
    transmit_buffer_1[227] = 8'h00;
    transmit_buffer_1[228] = 8'h00;
    transmit_buffer_1[229] = 8'h00;
    transmit_buffer_1[230] = 8'h00;
    transmit_buffer_1[231] = 8'h00;
    transmit_buffer_1[232] = 8'h00;
    transmit_buffer_1[233] = 8'h00;
    transmit_buffer_1[234] = 8'h00;
    transmit_buffer_1[235] = 8'h00;
    transmit_buffer_1[236] = 8'h00;
    transmit_buffer_1[237] = 8'h00;
    transmit_buffer_1[238] = 8'h00;
    transmit_buffer_1[239] = 8'h00;
    transmit_buffer_1[240] = 8'h00;
    transmit_buffer_1[241] = 8'h00;
    transmit_buffer_1[242] = 8'h00;
    transmit_buffer_1[243] = 8'h00;
    transmit_buffer_1[244] = 8'h00;
    transmit_buffer_1[245] = 8'h00;
    transmit_buffer_1[246] = 8'h00;
    transmit_buffer_1[247] = 8'h00;
    transmit_buffer_1[248] = 8'h00;
    transmit_buffer_1[249] = 8'h00;
    transmit_buffer_1[250] = 8'h00;
    transmit_buffer_1[251] = 8'h00;
    transmit_buffer_1[252] = 8'h00;
    transmit_buffer_1[253] = 8'h00;
    transmit_buffer_1[254] = 8'h00;
    transmit_buffer_1[255] = 8'h00;
    transmit_buffer_1[256] = 8'h00;
    transmit_buffer_1[257] = 8'h00;
    transmit_buffer_1[258] = 8'h00;
    transmit_buffer_1[259] = 8'h00;
    transmit_buffer_1[260] = 8'h00;
    transmit_buffer_1[261] = 8'h00;
    transmit_buffer_1[262] = 8'h00;
    transmit_buffer_1[263] = 8'h00;
    transmit_buffer_1[264] = 8'h00;
    transmit_buffer_1[265] = 8'h00;
    transmit_buffer_1[266] = 8'h00;
    transmit_buffer_1[267] = 8'h00;
    transmit_buffer_1[268] = 8'h00;
    transmit_buffer_1[269] = 8'h00;
    transmit_buffer_1[270] = 8'h00;
    transmit_buffer_1[271] = 8'h00;
    transmit_buffer_1[272] = 8'h00;
    transmit_buffer_1[273] = 8'h00;
    transmit_buffer_1[274] = 8'h00;
    transmit_buffer_1[275] = 8'h00;
    transmit_buffer_1[276] = 8'h00;
    transmit_buffer_1[277] = 8'h00;
    transmit_buffer_1[278] = 8'h00;
    transmit_buffer_1[279] = 8'h00;
    transmit_buffer_1[280] = 8'h00;
    transmit_buffer_1[281] = 8'h00;
    transmit_buffer_1[282] = 8'h00;
    transmit_buffer_1[283] = 8'h00;
    transmit_buffer_1[284] = 8'h00;
    transmit_buffer_1[285] = 8'h00;
    transmit_buffer_1[286] = 8'h00;
    transmit_buffer_1[287] = 8'h00;
    transmit_buffer_1[288] = 8'h00;
    transmit_buffer_1[289] = 8'h00;
    transmit_buffer_1[290] = 8'h00;
    transmit_buffer_1[291] = 8'h00;
    transmit_buffer_1[292] = 8'h00;
    transmit_buffer_1[293] = 8'h00;
    transmit_buffer_1[294] = 8'h00;
    transmit_buffer_1[295] = 8'h00;
    transmit_buffer_1[296] = 8'h00;
    transmit_buffer_1[297] = 8'h00;
    transmit_buffer_1[298] = 8'h00;
    transmit_buffer_1[299] = 8'h00;
    transmit_buffer_1[300] = 8'h00;
    transmit_buffer_1[301] = 8'h00;
    transmit_buffer_1[302] = 8'h00;
    transmit_buffer_1[303] = 8'h00;
    transmit_buffer_1[304] = 8'h00;
    transmit_buffer_1[305] = 8'h00;
    transmit_buffer_1[306] = 8'h00;
    transmit_buffer_1[307] = 8'h00;
    transmit_buffer_1[308] = 8'h00;
    transmit_buffer_1[309] = 8'h00;
    transmit_buffer_1[310] = 8'h00;
    transmit_buffer_1[311] = 8'h00;
    transmit_buffer_1[312] = 8'h00;
    transmit_buffer_1[313] = 8'h00;
    transmit_buffer_1[314] = 8'h00;
    transmit_buffer_1[315] = 8'h00;
    transmit_buffer_1[316] = 8'h00;
    transmit_buffer_1[317] = 8'h00;
    transmit_buffer_1[318] = 8'h00;
    transmit_buffer_1[319] = 8'h00;
    transmit_buffer_1[320] = 8'h00;
    transmit_buffer_1[321] = 8'h00;
    transmit_buffer_1[322] = 8'h00;
    transmit_buffer_1[323] = 8'h00;
    transmit_buffer_1[324] = 8'h00;
    transmit_buffer_1[325] = 8'h00;
    transmit_buffer_1[326] = 8'h00;
    transmit_buffer_1[327] = 8'h00;
    transmit_buffer_1[328] = 8'h00;
    transmit_buffer_1[329] = 8'h00;
    transmit_buffer_1[330] = 8'h00;
    transmit_buffer_1[331] = 8'h00;
    transmit_buffer_1[332] = 8'h00;
    transmit_buffer_1[333] = 8'h00;
    transmit_buffer_1[334] = 8'h00;
    transmit_buffer_1[335] = 8'h00;
    transmit_buffer_1[336] = 8'h00;
    transmit_buffer_1[337] = 8'h00;
    transmit_buffer_1[338] = 8'h00;
    transmit_buffer_1[339] = 8'h00;
    transmit_buffer_1[340] = 8'h00;
    transmit_buffer_1[341] = 8'h00;
    transmit_buffer_1[342] = 8'h00;
    transmit_buffer_1[343] = 8'h00;
    transmit_buffer_1[344] = 8'h00;
    transmit_buffer_1[345] = 8'h00;
    transmit_buffer_1[346] = 8'h00;
    transmit_buffer_1[347] = 8'h00;
    transmit_buffer_1[348] = 8'h00;
    transmit_buffer_1[349] = 8'h00;
    transmit_buffer_1[350] = 8'h00;
    transmit_buffer_1[351] = 8'h00;
    transmit_buffer_1[352] = 8'h00;
    transmit_buffer_1[353] = 8'h00;
    transmit_buffer_1[354] = 8'h00;
    transmit_buffer_1[355] = 8'h00;
    transmit_buffer_1[356] = 8'h00;
    transmit_buffer_1[357] = 8'h00;
    transmit_buffer_1[358] = 8'h00;
    transmit_buffer_1[359] = 8'h00;
    transmit_buffer_1[360] = 8'h00;
    transmit_buffer_1[361] = 8'h00;
    transmit_buffer_1[362] = 8'h00;
    transmit_buffer_1[363] = 8'h00;
    transmit_buffer_1[364] = 8'h00;
    transmit_buffer_1[365] = 8'h00;
    transmit_buffer_1[366] = 8'h00;
    transmit_buffer_1[367] = 8'h00;
    transmit_buffer_1[368] = 8'h00;
    transmit_buffer_1[369] = 8'h00;
    transmit_buffer_1[370] = 8'h00;
    transmit_buffer_1[371] = 8'h00;
    transmit_buffer_1[372] = 8'h00;
    transmit_buffer_1[373] = 8'h00;
    transmit_buffer_1[374] = 8'h00;
    transmit_buffer_1[375] = 8'h00;
    transmit_buffer_1[376] = 8'h00;
    transmit_buffer_1[377] = 8'h00;
    transmit_buffer_1[378] = 8'h00;
    transmit_buffer_1[379] = 8'h00;
    transmit_buffer_1[380] = 8'h00;
    transmit_buffer_1[381] = 8'h00;
    transmit_buffer_1[382] = 8'h00;
    transmit_buffer_1[383] = 8'h00;
    transmit_buffer_1[384] = 8'h00;
    transmit_buffer_1[385] = 8'h00;
    transmit_buffer_1[386] = 8'h00;
    transmit_buffer_1[387] = 8'h00;
    transmit_buffer_1[388] = 8'h00;
    transmit_buffer_1[389] = 8'h00;
    transmit_buffer_1[390] = 8'h00;
    transmit_buffer_1[391] = 8'h00;
    transmit_buffer_1[392] = 8'h00;
    transmit_buffer_1[393] = 8'h00;
    transmit_buffer_1[394] = 8'h00;
    transmit_buffer_1[395] = 8'h00;
    transmit_buffer_1[396] = 8'h00;
    transmit_buffer_1[397] = 8'h00;
    transmit_buffer_1[398] = 8'h00;
    transmit_buffer_1[399] = 8'h00;
    transmit_buffer_1[400] = 8'h00;
    transmit_buffer_1[401] = 8'h00;
    transmit_buffer_1[402] = 8'h00;
    transmit_buffer_1[403] = 8'h00;
    transmit_buffer_1[404] = 8'h00;
    transmit_buffer_1[405] = 8'h00;
    transmit_buffer_1[406] = 8'h00;
    transmit_buffer_1[407] = 8'h00;
    transmit_buffer_1[408] = 8'h00;
    transmit_buffer_1[409] = 8'h00;
    transmit_buffer_1[410] = 8'h00;
    transmit_buffer_1[411] = 8'h00;
    transmit_buffer_1[412] = 8'h00;
    transmit_buffer_1[413] = 8'h00;
    transmit_buffer_1[414] = 8'h00;
    transmit_buffer_1[415] = 8'h00;
    transmit_buffer_1[416] = 8'h00;
    transmit_buffer_1[417] = 8'h00;
    transmit_buffer_1[418] = 8'h00;
    transmit_buffer_1[419] = 8'h00;
    transmit_buffer_1[420] = 8'h00;
    transmit_buffer_1[421] = 8'h00;
    transmit_buffer_1[422] = 8'h00;
    transmit_buffer_1[423] = 8'h00;
    transmit_buffer_1[424] = 8'h00;
    transmit_buffer_1[425] = 8'h00;
    transmit_buffer_1[426] = 8'h00;
    transmit_buffer_1[427] = 8'h00;
    transmit_buffer_1[428] = 8'h00;
    transmit_buffer_1[429] = 8'h00;
    transmit_buffer_1[430] = 8'h00;
    transmit_buffer_1[431] = 8'h00;
    transmit_buffer_1[432] = 8'h00;
    transmit_buffer_1[433] = 8'h00;
    transmit_buffer_1[434] = 8'h00;
    transmit_buffer_1[435] = 8'h00;
    transmit_buffer_1[436] = 8'h00;
    transmit_buffer_1[437] = 8'h00;
    transmit_buffer_1[438] = 8'h00;
    transmit_buffer_1[439] = 8'h00;
    transmit_buffer_1[440] = 8'h00;
    transmit_buffer_1[441] = 8'h00;
    transmit_buffer_1[442] = 8'h00;
    transmit_buffer_1[443] = 8'h00;
    transmit_buffer_1[444] = 8'h00;
    transmit_buffer_1[445] = 8'h00;
    transmit_buffer_1[446] = 8'h00;
    transmit_buffer_1[447] = 8'h00;
    transmit_buffer_1[448] = 8'h00;
    transmit_buffer_1[449] = 8'h00;
    transmit_buffer_1[450] = 8'h00;
    transmit_buffer_1[451] = 8'h00;
    transmit_buffer_1[452] = 8'h00;
    transmit_buffer_1[453] = 8'h00;
    transmit_buffer_1[454] = 8'h00;
    transmit_buffer_1[455] = 8'h00;
    transmit_buffer_1[456] = 8'h00;
    transmit_buffer_1[457] = 8'h00;
    transmit_buffer_1[458] = 8'h00;
    transmit_buffer_1[459] = 8'h00;
    transmit_buffer_1[460] = 8'h00;
    transmit_buffer_1[461] = 8'h00;
    transmit_buffer_1[462] = 8'h00;
    transmit_buffer_1[463] = 8'h00;
    transmit_buffer_1[464] = 8'h00;
    transmit_buffer_1[465] = 8'h00;
    transmit_buffer_1[466] = 8'h00;
    transmit_buffer_1[467] = 8'h00;
    transmit_buffer_1[468] = 8'h00;
    transmit_buffer_1[469] = 8'h00;
    transmit_buffer_1[470] = 8'h00;
    transmit_buffer_1[471] = 8'h00;
    transmit_buffer_1[472] = 8'h00;
    transmit_buffer_1[473] = 8'h00;
    transmit_buffer_1[474] = 8'h00;
    transmit_buffer_1[475] = 8'h00;
    transmit_buffer_1[476] = 8'h00;
    transmit_buffer_1[477] = 8'h00;
    transmit_buffer_1[478] = 8'h00;
    transmit_buffer_1[479] = 8'h00;
    transmit_buffer_1[480] = 8'h00;
    transmit_buffer_1[481] = 8'h00;
    transmit_buffer_1[482] = 8'h00;
    transmit_buffer_1[483] = 8'h00;
    transmit_buffer_1[484] = 8'h00;
    transmit_buffer_1[485] = 8'h00;
    transmit_buffer_1[486] = 8'h00;
    transmit_buffer_1[487] = 8'h00;
    transmit_buffer_1[488] = 8'h00;
    transmit_buffer_1[489] = 8'h00;
    transmit_buffer_1[490] = 8'h00;
    transmit_buffer_1[491] = 8'h00;
    transmit_buffer_1[492] = 8'h00;
    transmit_buffer_1[493] = 8'h00;
    transmit_buffer_1[494] = 8'h00;
    transmit_buffer_1[495] = 8'h00;
    transmit_buffer_1[496] = 8'h00;
    transmit_buffer_1[497] = 8'h00;
    transmit_buffer_1[498] = 8'h00;
    transmit_buffer_1[499] = 8'h00;
    transmit_buffer_1[500] = 8'h00;
    transmit_buffer_1[501] = 8'h00;
    transmit_buffer_1[502] = 8'h00;
    transmit_buffer_1[503] = 8'h00;
    transmit_buffer_1[504] = 8'h00;
    transmit_buffer_1[505] = 8'h00;
    transmit_buffer_1[506] = 8'h00;
    transmit_buffer_1[507] = 8'h00;
    transmit_buffer_1[508] = 8'h00;
    transmit_buffer_1[509] = 8'h00;
    transmit_buffer_1[510] = 8'h00;
    transmit_buffer_1[511] = 8'h00;
  end
  always @(posedge usb_clk) begin
    if (transmit_buffer_1_w_en)
      transmit_buffer_1[transmit_buffer_1_w_addr] <= transmit_buffer_1_w_data;
  end
  reg [8:0] _1_;
  always @(posedge usb_clk) begin
    _1_ <= transmit_buffer_1_r_addr;
  end
  assign transmit_buffer_1_r_data = transmit_buffer_1[_1_];
  assign \$100  = generate_zlps &  \$98 ;
  assign \$102  = \$100  &  stream_ended_in_buffer1;
  assign \$104  = ~  ready;
  assign \$106  = \$signal$27  ==  10'h200;
  assign \$108  = generate_zlps &  \$106 ;
  assign \$110  = \$108  &  stream_ended_in_buffer1;
  assign \$112  = ~  ready;
  assign \$114  = \$signal  +  1'h1;
  assign \$116  = \$114  ==  10'h200;
  assign \$118  = \$116  |  last;
  assign \$11  = \$signal  +  1'h1;
  assign \$120  = valid &  \$118 ;
  assign \$122  = \$112  |  \$120 ;
  assign \$124  = ~  data_pid[0];
  assign \$126  = ~  data_pid[0];
  assign \$128  = \$signal$27  ==  10'h200;
  assign \$130  = generate_zlps &  \$128 ;
  assign \$132  = \$130  &  stream_ended_in_buffer1;
  assign \$134  = ~  ready;
  assign \$136  = \$signal$27  +  1'h1;
  assign \$138  = \$136  ==  10'h200;
  assign \$13  = \$11  ==  10'h200;
  assign \$140  = \$138  |  last;
  assign \$142  = valid &  \$140 ;
  assign \$144  = \$134  |  \$142 ;
  assign \$146  = ~  data_pid[0];
  assign \$148  = ~  data_pid[0];
  assign \$156  = ~  buffer_toggle;
  assign \$15  = \$13  |  last;
  assign \$159  = send_position +  1'h1;
  assign \$161  = ~  buffer_toggle;
  assign \$164  = send_position +  1'h1;
  assign \$167  = send_position +  1'h1;
  assign \$169  = ~  buffer_toggle;
  assign \$171  = \$signal  !=  10'h200;
  assign \$173  = ~  stream_ended_in_buffer0;
  assign \$175  = \$171  &  \$173 ;
  assign \$177  = \$signal$27  !=  10'h200;
  assign \$17  = valid &  \$15 ;
  assign \$179  = ~  stream_ended_in_buffer1;
  assign \$181  = \$177  &  \$179 ;
  assign \$183  = valid &  ready;
  assign \$185  = valid &  ready;
  assign \$187  = valid &  ready;
  assign \$190  = \$signal  +  1'h1;
  assign \$193  = \$signal$27  +  1'h1;
  assign \$195  = ~  buffer_toggle;
  assign \$197  = last &  transmit_buffer_0_w_en;
  assign \$19  = \$signal  +  1'h1;
  assign \$199  = last &  transmit_buffer_1_w_en;
  assign \$201  = \$signal  +  1'h1;
  assign \$203  = \$201  ==  10'h200;
  assign \$205  = \$203  |  last;
  assign \$207  = valid &  \$205 ;
  assign \$209  = \$signal  +  1'h1;
  assign \$211  = \$209  ==  10'h200;
  assign \$213  = \$211  |  last;
  assign \$217  = \$signal$27  +  1'h1;
  assign \$21  = \$19  ==  10'h200;
  assign \$219  = \$217  ==  10'h200;
  assign \$221  = \$219  |  last;
  assign \$223  = valid &  \$221 ;
  assign \$225  = \$signal$27  +  1'h1;
  assign \$227  = \$225  ==  10'h200;
  assign \$229  = \$227  |  last;
  assign \$233  = active &  is_in;
  assign \$235  = \$233  &  ready_for_response;
  assign \$238  = ~  buffer_toggle;
  assign \$23  = \$21  |  last;
  assign \$240  = |  \$signal ;
  assign \$242  = |  \$signal$27 ;
  assign \$244  = ~  buffer_toggle;
  assign \$246  = \$signal  ==  10'h200;
  assign \$248  = generate_zlps &  \$246 ;
  assign \$250  = \$248  &  stream_ended_in_buffer0;
  assign \$252  = ~  ready;
  assign \$254  = \$signal  ==  10'h200;
  assign \$256  = generate_zlps &  \$254 ;
  assign \$258  = \$256  &  stream_ended_in_buffer0;
  assign \$25  = ~  data_pid[0];
  assign \$260  = ~  ready;
  assign \$262  = \$signal  +  1'h1;
  assign \$264  = \$262  ==  10'h200;
  assign \$266  = \$264  |  last;
  assign \$268  = valid &  \$266 ;
  assign \$270  = \$260  |  \$268 ;
  assign \$272  = \$signal  ==  10'h200;
  assign \$274  = generate_zlps &  \$272 ;
  assign \$276  = \$274  &  stream_ended_in_buffer0;
  assign \$278  = ~  ready;
  assign \$280  = \$signal$27  +  1'h1;
  assign \$282  = \$280  ==  10'h200;
  assign \$284  = \$282  |  last;
  assign \$286  = valid &  \$284 ;
  assign \$288  = \$278  |  \$286 ;
  assign \$28  = \$signal$27  +  1'h1;
  assign \$290  = \$signal$27  ==  10'h200;
  assign \$292  = generate_zlps &  \$290 ;
  assign \$294  = \$292  &  stream_ended_in_buffer1;
  assign \$296  = ~  ready;
  assign \$298  = \$signal$27  ==  10'h200;
  assign \$300  = generate_zlps &  \$298 ;
  assign \$302  = \$300  &  stream_ended_in_buffer1;
  assign \$304  = ~  ready;
  assign \$306  = \$signal  +  1'h1;
  assign \$308  = \$306  ==  10'h200;
  assign \$30  = \$28  ==  10'h200;
  assign \$310  = \$308  |  last;
  assign \$312  = valid &  \$310 ;
  assign \$314  = \$304  |  \$312 ;
  assign \$316  = \$signal$27  ==  10'h200;
  assign \$318  = generate_zlps &  \$316 ;
  assign \$320  = \$318  &  stream_ended_in_buffer1;
  assign \$322  = ~  ready;
  assign \$324  = \$signal$27  +  1'h1;
  assign \$326  = \$324  ==  10'h200;
  assign \$328  = \$326  |  last;
  assign \$32  = \$30  |  last;
  assign \$330  = valid &  \$328 ;
  assign \$332  = \$322  |  \$330 ;
  assign \$334  = active &  is_in;
  assign \$336  = \$334  &  ready_for_response;
  assign \$338  = \$signal  +  1'h1;
  assign \$340  = \$338  ==  10'h200;
  assign \$342  = \$340  |  last;
  assign \$344  = valid &  \$342 ;
  assign \$346  = \$signal  +  1'h1;
  assign \$348  = \$346  ==  10'h200;
  assign \$34  = valid &  \$32 ;
  assign \$350  = \$348  |  last;
  assign \$352  = \$signal$27  +  1'h1;
  assign \$354  = \$352  ==  10'h200;
  assign \$356  = \$354  |  last;
  assign \$358  = valid &  \$356 ;
  assign \$360  = \$signal$27  +  1'h1;
  assign \$362  = \$360  ==  10'h200;
  assign \$364  = \$362  |  last;
  assign \$366  = active &  is_in;
  assign \$368  = \$366  &  ready_for_response;
  assign \$36  = \$signal$27  +  1'h1;
  assign \$371  = ~  buffer_toggle;
  assign \$373  = |  \$signal ;
  assign \$375  = |  \$signal$27 ;
  assign \$377  = send_position +  1'h1;
  assign \$379  = ~  buffer_toggle;
  assign \$381  = send_position +  1'h1;
  assign \$383  = \$381  ==  \$signal ;
  assign \$385  = send_position +  1'h1;
  assign \$387  = \$385  ==  \$signal$27 ;
  assign \$38  = \$36  ==  10'h200;
  assign \$389  = ~  buffer_toggle;
  assign \$391  = \$signal  ==  10'h200;
  assign \$393  = generate_zlps &  \$391 ;
  assign \$395  = \$393  &  stream_ended_in_buffer0;
  assign \$397  = ~  ready;
  assign \$399  = \$signal  ==  10'h200;
  assign \$401  = generate_zlps &  \$399 ;
  assign \$403  = \$401  &  stream_ended_in_buffer0;
  assign \$405  = ~  ready;
  assign \$407  = \$signal  +  1'h1;
  assign \$40  = \$38  |  last;
  assign \$409  = \$407  ==  10'h200;
  assign \$411  = \$409  |  last;
  assign \$413  = valid &  \$411 ;
  assign \$415  = \$405  |  \$413 ;
  assign \$417  = \$signal  ==  10'h200;
  assign \$419  = generate_zlps &  \$417 ;
  assign \$421  = \$419  &  stream_ended_in_buffer0;
  assign \$423  = ~  ready;
  assign \$425  = \$signal$27  +  1'h1;
  assign \$427  = \$425  ==  10'h200;
  assign \$42  = ~  data_pid[0];
  assign \$429  = \$427  |  last;
  assign \$431  = valid &  \$429 ;
  assign \$433  = \$423  |  \$431 ;
  assign \$435  = \$signal$27  ==  10'h200;
  assign \$437  = generate_zlps &  \$435 ;
  assign \$439  = \$437  &  stream_ended_in_buffer1;
  assign \$441  = ~  ready;
  assign \$443  = \$signal$27  ==  10'h200;
  assign \$445  = generate_zlps &  \$443 ;
  assign \$447  = \$445  &  stream_ended_in_buffer1;
  assign \$44  = ~  buffer_toggle;
  assign \$449  = ~  ready;
  assign \$451  = \$signal  +  1'h1;
  assign \$453  = \$451  ==  10'h200;
  assign \$455  = \$453  |  last;
  assign \$457  = valid &  \$455 ;
  assign \$459  = \$449  |  \$457 ;
  assign \$461  = \$signal$27  ==  10'h200;
  assign \$463  = generate_zlps &  \$461 ;
  assign \$465  = \$463  &  stream_ended_in_buffer1;
  assign \$467  = ~  ready;
  assign \$46  = \$signal  ==  10'h200;
  assign \$469  = \$signal$27  +  1'h1;
  assign \$471  = \$469  ==  10'h200;
  assign \$473  = \$471  |  last;
  assign \$475  = valid &  \$473 ;
  assign \$477  = \$467  |  \$475 ;
  assign \$479  = \$signal  +  1'h1;
  assign \$481  = \$479  ==  10'h200;
  assign \$483  = \$481  |  last;
  assign \$485  = valid &  \$483 ;
  assign \$487  = \$signal  +  1'h1;
  assign \$48  = generate_zlps &  \$46 ;
  assign \$489  = \$487  ==  10'h200;
  assign \$491  = \$489  |  last;
  assign \$495  = \$signal$27  +  1'h1;
  assign \$497  = \$495  ==  10'h200;
  assign \$499  = \$497  |  last;
  assign \$501  = valid &  \$499 ;
  assign \$503  = \$signal$27  +  1'h1;
  assign \$505  = \$503  ==  10'h200;
  assign \$507  = \$505  |  last;
  assign \$50  = \$48  &  stream_ended_in_buffer0;
  assign \$511  = ~  buffer_toggle;
  assign \$513  = \$signal  ==  10'h200;
  assign \$515  = generate_zlps &  \$513 ;
  assign \$517  = \$515  &  stream_ended_in_buffer0;
  assign \$519  = ~  ready;
  assign \$521  = \$signal  ==  10'h200;
  assign \$523  = generate_zlps &  \$521 ;
  assign \$525  = \$523  &  stream_ended_in_buffer0;
  assign \$527  = ~  ready;
  assign \$52  = ~  ready;
  assign \$529  = \$signal  +  1'h1;
  assign \$531  = \$529  ==  10'h200;
  assign \$533  = \$531  |  last;
  assign \$535  = valid &  \$533 ;
  assign \$537  = \$527  |  \$535 ;
  assign \$539  = \$signal  ==  10'h200;
  assign \$541  = generate_zlps &  \$539 ;
  assign \$543  = \$541  &  stream_ended_in_buffer0;
  assign \$545  = ~  ready;
  assign \$547  = \$signal$27  +  1'h1;
  assign \$54  = \$signal  ==  10'h200;
  assign \$549  = \$547  ==  10'h200;
  assign \$551  = \$549  |  last;
  assign \$553  = valid &  \$551 ;
  assign \$555  = \$545  |  \$553 ;
  assign \$557  = \$signal$27  ==  10'h200;
  assign \$559  = generate_zlps &  \$557 ;
  assign \$561  = \$559  &  stream_ended_in_buffer1;
  assign \$563  = ~  ready;
  assign \$565  = \$signal$27  ==  10'h200;
  assign \$567  = generate_zlps &  \$565 ;
  assign \$56  = generate_zlps &  \$54 ;
  assign \$569  = \$567  &  stream_ended_in_buffer1;
  assign \$571  = ~  ready;
  assign \$573  = \$signal  +  1'h1;
  assign \$575  = \$573  ==  10'h200;
  assign \$577  = \$575  |  last;
  assign \$579  = valid &  \$577 ;
  assign \$581  = \$571  |  \$579 ;
  assign \$583  = \$signal$27  ==  10'h200;
  assign \$585  = generate_zlps &  \$583 ;
  assign \$587  = \$585  &  stream_ended_in_buffer1;
  assign \$58  = \$56  &  stream_ended_in_buffer0;
  assign \$589  = ~  ready;
  assign \$591  = \$signal$27  +  1'h1;
  assign \$593  = \$591  ==  10'h200;
  assign \$595  = \$593  |  last;
  assign \$597  = valid &  \$595 ;
  assign \$599  = \$589  |  \$597 ;
  assign \$602  = send_position +  1'h1;
  assign \$604  = active &  is_in;
  assign \$606  = \$604  &  ready_for_response;
  assign \$60  = ~  ready;
  assign \$609  = ~  buffer_toggle;
  assign \$611  = |  \$signal ;
  assign \$613  = |  \$signal$27 ;
  assign \$615  = active &  is_in;
  assign \$617  = \$615  &  ready_for_response;
  assign \$620  = ~  buffer_toggle;
  assign \$622  = |  \$signal ;
  assign \$624  = |  \$signal$27 ;
  assign \$626  = active &  is_in;
  assign \$628  = \$626  &  ready_for_response;
  assign \$62  = \$signal  +  1'h1;
  assign \$631  = ~  buffer_toggle;
  assign \$633  = |  \$signal ;
  assign \$635  = |  \$signal$27 ;
  assign \$637  = send_position +  1'h1;
  assign \$639  = ~  buffer_toggle;
  assign \$641  = send_position +  1'h1;
  assign \$643  = \$641  ==  \$signal ;
  assign \$645  = send_position +  1'h1;
  assign \$647  = \$645  ==  \$signal$27 ;
  always @(posedge usb_clk)
    data_pid <= \data_pid$next ;
  assign \$64  = \$62  ==  10'h200;
  always @(posedge usb_clk)
    \$signal  <= \$signal$next ;
  always @(posedge usb_clk)
    \$signal$27  <= \$signal$27$next ;
  always @(posedge usb_clk)
    stream_ended_in_buffer0 <= \stream_ended_in_buffer0$next ;
  always @(posedge usb_clk)
    stream_ended_in_buffer1 <= \stream_ended_in_buffer1$next ;
  always @(posedge usb_clk)
    fsm_state <= \fsm_state$next ;
  always @(posedge usb_clk)
    buffer_toggle <= \buffer_toggle$next ;
  always @(posedge usb_clk)
    send_position <= \send_position$next ;
  always @(posedge usb_clk)
    first <= \first$next ;
  assign \$66  = \$64  |  last;
  assign \$68  = valid &  \$66 ;
  assign \$70  = \$60  |  \$68 ;
  assign \$72  = ~  data_pid[0];
  assign \$74  = ~  data_pid[0];
  assign \$76  = \$signal  ==  10'h200;
  assign \$78  = generate_zlps &  \$76 ;
  assign \$80  = \$78  &  stream_ended_in_buffer0;
  assign \$82  = ~  ready;
  assign \$84  = \$signal$27  +  1'h1;
  assign \$86  = \$84  ==  10'h200;
  assign \$88  = \$86  |  last;
  assign \$90  = valid &  \$88 ;
  assign \$92  = \$82  |  \$90 ;
  assign \$94  = ~  data_pid[0];
  assign \$96  = ~  data_pid[0];
  assign \$98  = \$signal$27  ==  10'h200;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$32 ) begin end
    \data_pid$next  = data_pid;
    casez (reset_sequence)
      1'h1:
          \data_pid$next  = \$7 ;
    endcase
    casez (fsm_state)
      2'h0:
          casez (buffer_toggle)
            1'h0:
                casez (\$17 )
                  1'h1:
                      casez (\$23 )
                        1'h1:
                            \data_pid$next [0] = \$25 ;
                      endcase
                endcase
            1'h?:
                casez (\$34 )
                  1'h1:
                      casez (\$40 )
                        1'h1:
                            \data_pid$next [0] = \$42 ;
                      endcase
                endcase
          endcase
      2'h1:
          ;
      2'h2:
          ;
      2'h3:
          casez (ack)
            1'h1:
                casez (\$44 )
                  1'h0:
                      casez (buffer_toggle)
                        1'h0:
                            casez ({ \$70 , \$58  })
                              2'b?1:
                                  \data_pid$next [0] = \$72 ;
                              2'b1?:
                                  \data_pid$next [0] = \$74 ;
                            endcase
                        1'h?:
                            casez ({ \$92 , \$80  })
                              2'b?1:
                                  \data_pid$next [0] = \$94 ;
                              2'b1?:
                                  \data_pid$next [0] = \$96 ;
                            endcase
                      endcase
                  1'h?:
                      casez (buffer_toggle)
                        1'h0:
                            casez ({ \$122 , \$110  })
                              2'b?1:
                                  \data_pid$next [0] = \$124 ;
                              2'b1?:
                                  \data_pid$next [0] = \$126 ;
                            endcase
                        1'h?:
                            casez ({ \$144 , \$132  })
                              2'b?1:
                                  \data_pid$next [0] = \$146 ;
                              2'b1?:
                                  \data_pid$next [0] = \$148 ;
                            endcase
                      endcase
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \data_pid$next  = 2'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$32 ) begin end
    \$signal$next  = \$signal ;
    \$signal$27$next  = \$signal$27 ;
    casez (buffer_toggle)
      1'h0:
          casez (transmit_buffer_0_w_en)
            1'h1:
                \$signal$next  = \$190 [9:0];
          endcase
      1'h?:
          casez (transmit_buffer_1_w_en)
            1'h1:
                \$signal$27$next  = \$193 [9:0];
          endcase
    endcase
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          ;
      2'h2:
          ;
      2'h3:
          casez (ack)
            1'h1:
                casez (\$195 )
                  1'h0:
                      \$signal$next  = 10'h000;
                  1'h?:
                      \$signal$27$next  = 10'h000;
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
        begin
          \$signal$next  = 10'h000;
          \$signal$27$next  = 10'h000;
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$32 ) begin end
    \stream_ended_in_buffer0$next  = stream_ended_in_buffer0;
    \stream_ended_in_buffer1$next  = stream_ended_in_buffer1;
    casez (buffer_toggle)
      1'h0:
          casez (\$197 )
            1'h1:
                \stream_ended_in_buffer0$next  = 1'h1;
          endcase
      1'h?:
          casez (\$199 )
            1'h1:
                \stream_ended_in_buffer1$next  = 1'h1;
          endcase
    endcase
    casez (fsm_state)
      2'h0:
          casez (buffer_toggle)
            1'h0:
                casez (\$207 )
                  1'h1:
                      casez (\$213 )
                        1'h1:
                            casez (\$215 )
                              1'h0:
                                  \stream_ended_in_buffer0$next  = 1'h0;
                              1'h?:
                                  \stream_ended_in_buffer1$next  = 1'h0;
                            endcase
                      endcase
                endcase
            1'h?:
                casez (\$223 )
                  1'h1:
                      casez (\$229 )
                        1'h1:
                            casez (\$231 )
                              1'h0:
                                  \stream_ended_in_buffer0$next  = 1'h0;
                              1'h?:
                                  \stream_ended_in_buffer1$next  = 1'h0;
                            endcase
                      endcase
                endcase
          endcase
      2'h1:
          casez (\$235 )
            1'h1:
                casez (\$238 )
                  1'h0:
                      casez (\$240 )
                        1'h1:
                            ;
                        default:
                            \stream_ended_in_buffer0$next  = 1'h0;
                      endcase
                  1'h?:
                      casez (\$242 )
                        1'h1:
                            ;
                        default:
                            \stream_ended_in_buffer1$next  = 1'h0;
                      endcase
                endcase
          endcase
      2'h2:
          ;
      2'h3:
          casez (ack)
            1'h1:
                casez (\$244 )
                  1'h0:
                      casez (buffer_toggle)
                        1'h0:
                            casez ({ \$270 , \$258  })
                              2'b?1:
                                  ;
                              2'b1?:
                                  \stream_ended_in_buffer0$next  = 1'h0;
                            endcase
                        1'h?:
                            casez ({ \$288 , \$276  })
                              2'b?1:
                                  ;
                              2'b1?:
                                  \stream_ended_in_buffer0$next  = 1'h0;
                            endcase
                      endcase
                  1'h?:
                      casez (buffer_toggle)
                        1'h0:
                            casez ({ \$314 , \$302  })
                              2'b?1:
                                  ;
                              2'b1?:
                                  \stream_ended_in_buffer1$next  = 1'h0;
                            endcase
                        1'h?:
                            casez ({ \$332 , \$320  })
                              2'b?1:
                                  ;
                              2'b1?:
                                  \stream_ended_in_buffer1$next  = 1'h0;
                            endcase
                      endcase
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
        begin
          \stream_ended_in_buffer0$next  = 1'h0;
          \stream_ended_in_buffer1$next  = 1'h0;
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$32 ) begin end
    nak = 1'h0;
    casez (fsm_state)
      2'h0:
          nak = \$336 ;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$32 ) begin end
    \fsm_state$next  = fsm_state;
    casez (fsm_state)
      2'h0:
          casez (buffer_toggle)
            1'h0:
                casez (\$344 )
                  1'h1:
                      casez (\$350 )
                        1'h1:
                            \fsm_state$next  = 2'h1;
                      endcase
                endcase
            1'h?:
                casez (\$358 )
                  1'h1:
                      casez (\$364 )
                        1'h1:
                            \fsm_state$next  = 2'h1;
                      endcase
                endcase
          endcase
      2'h1:
          casez (\$368 )
            1'h1:
                casez (\$371 )
                  1'h0:
                      casez (\$373 )
                        1'h1:
                            \fsm_state$next  = 2'h2;
                        default:
                            \fsm_state$next  = 2'h3;
                      endcase
                  1'h?:
                      casez (\$375 )
                        1'h1:
                            \fsm_state$next  = 2'h2;
                        default:
                            \fsm_state$next  = 2'h3;
                      endcase
                endcase
          endcase
      2'h2:
          casez (\ready$4 )
            1'h1:
                casez (\$379 )
                  1'h0:
                      casez (\$383 )
                        1'h1:
                            \fsm_state$next  = 2'h3;
                      endcase
                  1'h?:
                      casez (\$387 )
                        1'h1:
                            \fsm_state$next  = 2'h3;
                      endcase
                endcase
          endcase
      2'h3:
        begin
          casez (ack)
            1'h1:
                casez (\$389 )
                  1'h0:
                      casez (buffer_toggle)
                        1'h0:
                            casez ({ \$415 , \$403  })
                              2'b?1:
                                  \fsm_state$next  = 2'h1;
                              2'b1?:
                                  \fsm_state$next  = 2'h1;
                              default:
                                  \fsm_state$next  = 2'h0;
                            endcase
                        1'h?:
                            casez ({ \$433 , \$421  })
                              2'b?1:
                                  \fsm_state$next  = 2'h1;
                              2'b1?:
                                  \fsm_state$next  = 2'h1;
                              default:
                                  \fsm_state$next  = 2'h0;
                            endcase
                      endcase
                  1'h?:
                      casez (buffer_toggle)
                        1'h0:
                            casez ({ \$459 , \$447  })
                              2'b?1:
                                  \fsm_state$next  = 2'h1;
                              2'b1?:
                                  \fsm_state$next  = 2'h1;
                              default:
                                  \fsm_state$next  = 2'h0;
                            endcase
                        1'h?:
                            casez ({ \$477 , \$465  })
                              2'b?1:
                                  \fsm_state$next  = 2'h1;
                              2'b1?:
                                  \fsm_state$next  = 2'h1;
                              default:
                                  \fsm_state$next  = 2'h0;
                            endcase
                      endcase
                endcase
          endcase
          casez (new_token)
            1'h1:
                \fsm_state$next  = 2'h1;
          endcase
        end
    endcase
    casez (usb_rst)
      1'h1:
          \fsm_state$next  = 2'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$32 ) begin end
    \buffer_toggle$next  = buffer_toggle;
    casez (fsm_state)
      2'h0:
          casez (buffer_toggle)
            1'h0:
                casez (\$485 )
                  1'h1:
                      casez (\$491 )
                        1'h1:
                            \buffer_toggle$next  = \$493 ;
                      endcase
                endcase
            1'h?:
                casez (\$501 )
                  1'h1:
                      casez (\$507 )
                        1'h1:
                            \buffer_toggle$next  = \$509 ;
                      endcase
                endcase
          endcase
      2'h1:
          ;
      2'h2:
          ;
      2'h3:
          casez (ack)
            1'h1:
                casez (\$511 )
                  1'h0:
                      casez (buffer_toggle)
                        1'h0:
                            casez ({ \$537 , \$525  })
                              2'b?1:
                                  ;
                              2'b1?:
                                  \buffer_toggle$next  = 1'h0;
                            endcase
                        1'h?:
                            casez ({ \$555 , \$543  })
                              2'b?1:
                                  ;
                              2'b1?:
                                  \buffer_toggle$next  = 1'h0;
                            endcase
                      endcase
                  1'h?:
                      casez (buffer_toggle)
                        1'h0:
                            casez ({ \$581 , \$569  })
                              2'b?1:
                                  ;
                              2'b1?:
                                  \buffer_toggle$next  = 1'h1;
                            endcase
                        1'h?:
                            casez ({ \$599 , \$587  })
                              2'b?1:
                                  ;
                              2'b1?:
                                  \buffer_toggle$next  = 1'h1;
                            endcase
                      endcase
                endcase
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \buffer_toggle$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$32 ) begin end
    \send_position$next  = send_position;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          \send_position$next  = 10'h000;
      2'h2:
          casez (\ready$4 )
            1'h1:
                \send_position$next  = \$602 [9:0];
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \send_position$next  = 10'h000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$32 ) begin end
    \first$next  = first;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          casez (\$606 )
            1'h1:
                casez (\$609 )
                  1'h0:
                      casez (\$611 )
                        1'h1:
                            \first$next  = 1'h1;
                      endcase
                  1'h?:
                      casez (\$613 )
                        1'h1:
                            \first$next  = 1'h1;
                      endcase
                endcase
          endcase
      2'h2:
          casez (\ready$4 )
            1'h1:
                \first$next  = 1'h0;
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \first$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$32 ) begin end
    casez (buffer_toggle)
      1'h0:
          transmit_buffer_0_w_addr = \$signal [8:0];
      1'h?:
          transmit_buffer_0_w_addr = \$signal$27 [8:0];
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$32 ) begin end
    \valid$1  = 1'h0;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          casez (\$617 )
            1'h1:
                casez (\$620 )
                  1'h0:
                      casez (\$622 )
                        1'h1:
                            ;
                        default:
                            \valid$1  = 1'h1;
                      endcase
                  1'h?:
                      casez (\$624 )
                        1'h1:
                            ;
                        default:
                            \valid$1  = 1'h1;
                      endcase
                endcase
          endcase
      2'h2:
          \valid$1  = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$32 ) begin end
    \last$2  = 1'h0;
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          casez (\$628 )
            1'h1:
                casez (\$631 )
                  1'h0:
                      casez (\$633 )
                        1'h1:
                            ;
                        default:
                            \last$2  = 1'h1;
                      endcase
                  1'h?:
                      casez (\$635 )
                        1'h1:
                            ;
                        default:
                            \last$2  = 1'h1;
                      endcase
                endcase
          endcase
      2'h2:
          casez (\$639 )
            1'h0:
                \last$2  = \$643 ;
            1'h?:
                \last$2  = \$647 ;
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$32 ) begin end
    casez (buffer_toggle)
      1'h0:
          transmit_buffer_1_w_addr = \$signal [8:0];
      1'h?:
          transmit_buffer_1_w_addr = \$signal$27 [8:0];
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$32 ) begin end
    transmit_buffer_0_r_addr = 9'h000;
    transmit_buffer_1_r_addr = 9'h000;
    casez (\$156 )
      1'h0:
          transmit_buffer_0_r_addr = send_position[8:0];
      1'h?:
          transmit_buffer_1_r_addr = send_position[8:0];
    endcase
    casez (fsm_state)
      2'h0:
          ;
      2'h1:
          ;
      2'h2:
          casez (\ready$4 )
            1'h1:
                casez (\$161 )
                  1'h0:
                      transmit_buffer_0_r_addr = \$164 [8:0];
                  1'h?:
                      transmit_buffer_1_r_addr = \$167 [8:0];
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$32 ) begin end
    casez (\$169 )
      1'h0:
          \payload$3  = transmit_buffer_0_r_data;
      1'h?:
          \payload$3  = transmit_buffer_1_r_data;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$32 ) begin end
    casez (buffer_toggle)
      1'h0:
          ready = \$175 ;
      1'h?:
          ready = \$181 ;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$32 ) begin end
    transmit_buffer_0_w_en = 1'h0;
    transmit_buffer_1_w_en = 1'h0;
    casez (buffer_toggle)
      1'h0:
          transmit_buffer_0_w_en = \$185 ;
      1'h?:
          transmit_buffer_1_w_en = \$187 ;
    endcase
  end
  assign \$151  = \$signal ;
  assign \$152  = \$signal$27 ;
  assign \$154  = \$signal ;
  assign \$155  = \$signal$27 ;
  assign \$158  = \$159 ;
  assign \$163  = \$164 ;
  assign \$166  = \$167 ;
  assign \$189  = \$190 ;
  assign \$192  = \$193 ;
  assign \$601  = \$602 ;
  assign reset_sequence = 1'h0;
  assign start_with_data1 = 1'h0;
  assign transmit_buffer_1_w_data = payload;
  assign transmit_buffer_0_w_data = payload;
  assign \$8  = 1'h1;
  assign \$7  = 2'h1;
  assign \$215  = 1'h1;
  assign \$231  = 1'h0;
  assign \$493  = 1'h1;
  assign \$509  = 1'h0;
endmodule
module tx_multiplexer(valid, ready, \valid$1 , \data$2 , \data$3 , \valid$4 , \ready$5 , \valid$6 , \data$7 , \ready$8 , data);
  reg \$auto$verilog_backend.cc:2083:dump_module$33  = 0;
  wire \$11 ;
  wire \$13 ;
  wire \$9 ;
  output [7:0] data;
  reg [7:0] data;
  input [7:0] \data$2 ;
  wire [7:0] \data$2 ;
  input [7:0] \data$3 ;
  wire [7:0] \data$3 ;
  input [7:0] \data$7 ;
  wire [7:0] \data$7 ;
  wire [2:0] encoder_i;
  wire [1:0] encoder_o;
  input ready;
  wire ready;
  wire \ready$15 ;
  output \ready$5 ;
  wire \ready$5 ;
  output \ready$8 ;
  wire \ready$8 ;
  output valid;
  wire valid;
  input \valid$1 ;
  wire \valid$1 ;
  input \valid$4 ;
  wire \valid$4 ;
  input \valid$6 ;
  wire \valid$6 ;
  assign \$11  = \$9  |  \valid$4 ;
  assign \$13  = \$11  |  \valid$6 ;
  \encoder$6  encoder (
    .i(encoder_i),
    .o(encoder_o)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$33 ) begin end
    data = 8'h00;
    casez (encoder_o)
      2'h0:
          data = \data$2 ;
      2'h1:
          data = \data$3 ;
      2'h2:
          data = \data$7 ;
    endcase
  end
  assign \ready$8  = ready;
  assign \ready$5  = ready;
  assign \ready$15  = ready;
  assign valid = \$13 ;
  assign encoder_i[2] = \valid$6 ;
  assign encoder_i[1] = \valid$4 ;
  assign encoder_i[0] = \valid$1 ;
  assign \$9  = \valid$1 ;
endmodule
module tx_mux(first, last, payload, ready, \valid$1 , \valid$2 , \valid$3 , \valid$4 , \payload$5 , \payload$6 , \payload$7 , \first$8 , \first$9 , \first$10 , \last$11 , \last$12 , \last$13 , \ready$14 , \ready$15 , \ready$16 , valid
);
  reg \$auto$verilog_backend.cc:2083:dump_module$34  = 0;
  wire \$18 ;
  wire \$20 ;
  wire \$22 ;
  wire \$24 ;
  wire \$26 ;
  wire \$28 ;
  wire \$31 ;
  wire \$33 ;
  wire \$35 ;
  wire \$37 ;
  wire \$40 ;
  wire \$42 ;
  wire [3:0] encoder_i;
  wire [1:0] encoder_o;
  output first;
  wire first;
  input \first$10 ;
  wire \first$10 ;
  wire \first$30 ;
  input \first$8 ;
  wire \first$8 ;
  input \first$9 ;
  wire \first$9 ;
  output last;
  wire last;
  input \last$11 ;
  wire \last$11 ;
  input \last$12 ;
  wire \last$12 ;
  input \last$13 ;
  wire \last$13 ;
  wire \last$39 ;
  output [7:0] payload;
  reg [7:0] payload;
  wire [7:0] \payload$17 ;
  input [7:0] \payload$5 ;
  wire [7:0] \payload$5 ;
  input [7:0] \payload$6 ;
  wire [7:0] \payload$6 ;
  input [7:0] \payload$7 ;
  wire [7:0] \payload$7 ;
  input ready;
  wire ready;
  output \ready$14 ;
  wire \ready$14 ;
  output \ready$15 ;
  wire \ready$15 ;
  output \ready$16 ;
  wire \ready$16 ;
  wire \ready$44 ;
  output valid;
  wire valid;
  input \valid$1 ;
  wire \valid$1 ;
  input \valid$2 ;
  wire \valid$2 ;
  input \valid$3 ;
  wire \valid$3 ;
  input \valid$4 ;
  wire \valid$4 ;
  assign \$20  = \$18  |  \valid$2 ;
  assign \$22  = \$20  |  \valid$3 ;
  assign \$24  = \$22  |  \valid$4 ;
  assign \$28  = \$26  |  \first$9 ;
  assign \$33  = \$31  |  \first$10 ;
  assign \$37  = \$35  |  \last$12 ;
  assign \$42  = \$40  |  \last$13 ;
  encoder encoder (
    .i(encoder_i),
    .o(encoder_o)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$34 ) begin end
    casez (encoder_o)
      2'h0:
          payload = \payload$5 ;
      2'h1:
          payload = \payload$6 ;
      2'h2:
          payload = 8'h00;
      2'h3:
          payload = \payload$7 ;
    endcase
  end
  assign \payload$17  = 8'h00;
  assign \first$30  = 1'h0;
  assign \last$39  = 1'h0;
  assign \ready$16  = ready;
  assign \ready$44  = ready;
  assign \ready$15  = ready;
  assign \ready$14  = ready;
  assign last = \$42 ;
  assign first = \$33 ;
  assign valid = \$24 ;
  assign encoder_i[3] = \valid$4 ;
  assign encoder_i[2] = \valid$3 ;
  assign encoder_i[1] = \valid$2 ;
  assign encoder_i[0] = \valid$1 ;
  assign \$18  = \valid$1 ;
  assign \$26  = \first$8 ;
  assign \$31  = \$28 ;
  assign \$35  = \last$11 ;
  assign \$40  = \$37 ;
endmodule
module \tx_mux$2 (first, last, payload, ready, \valid$1 , \valid$2 , \valid$3 , \payload$4 , \first$5 , \last$6 , \last$7 , \ready$8 , valid);
  reg \$auto$verilog_backend.cc:2083:dump_module$35  = 0;
  wire \$11 ;
  wire \$13 ;
  wire \$15 ;
  wire \$17 ;
  wire \$20 ;
  wire \$23 ;
  wire \$25 ;
  wire \$27 ;
  wire \$30 ;
  wire [2:0] encoder_i;
  wire [1:0] encoder_o;
  output first;
  wire first;
  wire \first$19 ;
  wire \first$22 ;
  input \first$5 ;
  wire \first$5 ;
  output last;
  wire last;
  wire \last$29 ;
  input \last$6 ;
  wire \last$6 ;
  input \last$7 ;
  wire \last$7 ;
  output [7:0] payload;
  reg [7:0] payload;
  wire [7:0] \payload$10 ;
  input [7:0] \payload$4 ;
  wire [7:0] \payload$4 ;
  wire [7:0] \payload$9 ;
  input ready;
  wire ready;
  wire \ready$32 ;
  wire \ready$33 ;
  output \ready$8 ;
  wire \ready$8 ;
  output valid;
  wire valid;
  input \valid$1 ;
  wire \valid$1 ;
  input \valid$2 ;
  wire \valid$2 ;
  input \valid$3 ;
  wire \valid$3 ;
  assign \$13  = \$11  |  \valid$2 ;
  assign \$15  = \$13  |  \valid$3 ;
  assign \$27  = \$25  |  \last$7 ;
  \encoder$3  encoder (
    .i(encoder_i),
    .o(encoder_o)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$35 ) begin end
    payload = 8'h00;
    casez (encoder_o)
      2'h0:
          payload = \payload$4 ;
      2'h1:
          payload = 8'h00;
      2'h2:
          payload = 8'h00;
    endcase
  end
  assign \payload$9  = 8'h00;
  assign \payload$10  = 8'h00;
  assign \first$19  = 1'h0;
  assign \first$22  = 1'h0;
  assign \last$29  = 1'h0;
  assign \ready$33  = ready;
  assign \ready$32  = ready;
  assign \ready$8  = ready;
  assign last = \$30 ;
  assign first = \$23 ;
  assign valid = \$15 ;
  assign encoder_i[2] = \valid$3 ;
  assign encoder_i[1] = \valid$2 ;
  assign encoder_i[0] = \valid$1 ;
  assign \$11  = \valid$1 ;
  assign \$17  = \first$5 ;
  assign \$20  = \first$5 ;
  assign \$23  = \first$5 ;
  assign \$25  = \last$6 ;
  assign \$30  = \$27 ;
endmodule
module usb(first, last, payload, ready, \valid$1 , \first$2 , \last$3 , \payload$4 , \ready$5 , connect, usb_rst, usb_clk, ulpi__clk, ulpi__rst, ulpi__data__oe, ulpi__dir__i, ulpi__nxt, ulpi__data__i, ulpi__data__o, ulpi__stp, valid
);
  reg \$auto$verilog_backend.cc:2083:dump_module$36  = 0;
  wire \$111 ;
  wire [1:0] \$113 ;
  wire \$115 ;
  wire [1:0] \$117 ;
  wire [1:0] \$118 ;
  wire [1:0] \$120 ;
  wire \$122 ;
  wire \$124 ;
  wire \$126 ;
  wire [3:0] \$128 ;
  wire [3:0] \$129 ;
  reg [6:0] address = 7'h00;
  reg [6:0] \address$next ;
  reg [7:0] configuration = 8'h00;
  reg [7:0] \configuration$next ;
  input connect;
  wire connect;
  wire [15:0] data_crc_crc;
  wire [7:0] data_crc_rx_data;
  wire data_crc_rx_valid;
  wire data_crc_start;
  wire [7:0] data_crc_tx_data;
  wire data_crc_tx_valid;
  wire endpoint_mux_ack;
  wire \endpoint_mux_ack$12 ;
  wire \endpoint_mux_ack$15 ;
  wire \endpoint_mux_ack$36 ;
  wire \endpoint_mux_ack$62 ;
  wire \endpoint_mux_ack$81 ;
  wire \endpoint_mux_ack$82 ;
  wire \endpoint_mux_ack$83 ;
  wire \endpoint_mux_ack$84 ;
  wire [6:0] endpoint_mux_active_address;
  wire [7:0] endpoint_mux_active_config;
  wire [7:0] \endpoint_mux_active_config$35 ;
  wire [6:0] endpoint_mux_address;
  wire [6:0] \endpoint_mux_address$20 ;
  wire [6:0] \endpoint_mux_address$41 ;
  wire [6:0] \endpoint_mux_address$67 ;
  wire endpoint_mux_address_changed;
  wire \endpoint_mux_address_changed$77 ;
  wire endpoint_mux_config_changed;
  wire \endpoint_mux_config_changed$79 ;
  wire [15:0] endpoint_mux_crc;
  wire [3:0] endpoint_mux_endpoint;
  wire [3:0] \endpoint_mux_endpoint$21 ;
  wire [3:0] \endpoint_mux_endpoint$42 ;
  wire [3:0] \endpoint_mux_endpoint$51 ;
  wire [3:0] \endpoint_mux_endpoint$68 ;
  wire endpoint_mux_first;
  wire \endpoint_mux_first$102 ;
  wire \endpoint_mux_first$103 ;
  wire \endpoint_mux_first$104 ;
  wire [10:0] endpoint_mux_frame;
  wire [10:0] \endpoint_mux_frame$24 ;
  wire [10:0] \endpoint_mux_frame$45 ;
  wire [10:0] \endpoint_mux_frame$71 ;
  wire endpoint_mux_is_in;
  wire \endpoint_mux_is_in$26 ;
  wire \endpoint_mux_is_in$47 ;
  wire \endpoint_mux_is_in$73 ;
  wire endpoint_mux_is_out;
  wire \endpoint_mux_is_out$27 ;
  wire \endpoint_mux_is_out$48 ;
  wire \endpoint_mux_is_out$53 ;
  wire \endpoint_mux_is_out$74 ;
  wire endpoint_mux_is_ping;
  wire \endpoint_mux_is_ping$29 ;
  wire \endpoint_mux_is_ping$50 ;
  wire \endpoint_mux_is_ping$54 ;
  wire \endpoint_mux_is_ping$76 ;
  wire endpoint_mux_is_setup;
  wire \endpoint_mux_is_setup$28 ;
  wire \endpoint_mux_is_setup$49 ;
  wire \endpoint_mux_is_setup$75 ;
  wire endpoint_mux_last;
  wire \endpoint_mux_last$105 ;
  wire \endpoint_mux_last$106 ;
  wire \endpoint_mux_last$107 ;
  wire endpoint_mux_nak;
  wire \endpoint_mux_nak$13 ;
  wire \endpoint_mux_nak$16 ;
  wire \endpoint_mux_nak$37 ;
  wire \endpoint_mux_nak$63 ;
  wire \endpoint_mux_nak$85 ;
  wire \endpoint_mux_nak$86 ;
  wire \endpoint_mux_nak$87 ;
  wire \endpoint_mux_nak$88 ;
  wire [6:0] endpoint_mux_new_address;
  wire [6:0] \endpoint_mux_new_address$78 ;
  wire [7:0] endpoint_mux_new_config;
  wire [7:0] \endpoint_mux_new_config$80 ;
  wire endpoint_mux_new_frame;
  wire \endpoint_mux_new_frame$25 ;
  wire \endpoint_mux_new_frame$46 ;
  wire \endpoint_mux_new_frame$72 ;
  wire endpoint_mux_new_token;
  wire \endpoint_mux_new_token$22 ;
  wire \endpoint_mux_new_token$43 ;
  wire \endpoint_mux_new_token$69 ;
  wire endpoint_mux_next;
  wire \endpoint_mux_next$31 ;
  wire \endpoint_mux_next$56 ;
  wire endpoint_mux_nyet;
  wire \endpoint_mux_nyet$18 ;
  wire \endpoint_mux_nyet$39 ;
  wire \endpoint_mux_nyet$65 ;
  wire [7:0] endpoint_mux_payload;
  wire [7:0] \endpoint_mux_payload$100 ;
  wire [7:0] \endpoint_mux_payload$101 ;
  wire [7:0] \endpoint_mux_payload$11 ;
  wire [7:0] \endpoint_mux_payload$32 ;
  wire [7:0] \endpoint_mux_payload$57 ;
  wire [7:0] \endpoint_mux_payload$99 ;
  wire [3:0] endpoint_mux_pid;
  wire [3:0] \endpoint_mux_pid$19 ;
  wire [3:0] \endpoint_mux_pid$40 ;
  wire [3:0] \endpoint_mux_pid$66 ;
  wire endpoint_mux_ready;
  wire \endpoint_mux_ready$108 ;
  wire \endpoint_mux_ready$109 ;
  wire \endpoint_mux_ready$110 ;
  wire endpoint_mux_ready_for_response;
  wire \endpoint_mux_ready_for_response$23 ;
  wire \endpoint_mux_ready_for_response$44 ;
  wire \endpoint_mux_ready_for_response$52 ;
  wire \endpoint_mux_ready_for_response$70 ;
  wire endpoint_mux_rx_complete;
  wire \endpoint_mux_rx_complete$58 ;
  wire endpoint_mux_rx_invalid;
  wire \endpoint_mux_rx_invalid$60 ;
  wire [1:0] endpoint_mux_rx_pid_toggle;
  wire [1:0] \endpoint_mux_rx_pid_toggle$61 ;
  wire endpoint_mux_rx_ready_for_response;
  wire \endpoint_mux_rx_ready_for_response$33 ;
  wire \endpoint_mux_rx_ready_for_response$59 ;
  wire endpoint_mux_rx_timeout;
  wire [1:0] endpoint_mux_speed;
  wire [1:0] \endpoint_mux_speed$34 ;
  wire endpoint_mux_stall;
  wire \endpoint_mux_stall$14 ;
  wire \endpoint_mux_stall$17 ;
  wire \endpoint_mux_stall$38 ;
  wire \endpoint_mux_stall$64 ;
  wire \endpoint_mux_stall$89 ;
  wire \endpoint_mux_stall$90 ;
  wire \endpoint_mux_stall$91 ;
  wire endpoint_mux_start;
  wire \endpoint_mux_start$92 ;
  wire endpoint_mux_tx_allowed;
  wire [1:0] endpoint_mux_tx_pid_toggle;
  wire [1:0] \endpoint_mux_tx_pid_toggle$96 ;
  wire [1:0] \endpoint_mux_tx_pid_toggle$97 ;
  wire [1:0] \endpoint_mux_tx_pid_toggle$98 ;
  wire endpoint_mux_tx_timeout;
  wire endpoint_mux_valid;
  wire \endpoint_mux_valid$10 ;
  wire \endpoint_mux_valid$30 ;
  wire \endpoint_mux_valid$55 ;
  wire \endpoint_mux_valid$93 ;
  wire \endpoint_mux_valid$94 ;
  wire \endpoint_mux_valid$95 ;
  input first;
  wire first;
  output \first$2 ;
  wire \first$2 ;
  reg [10:0] frame_number = 11'h000;
  reg [10:0] \frame_number$next ;
  wire full_speed_only;
  wire handshake_detector_ack;
  wire handshake_detector_nak;
  wire handshake_detector_nyet;
  wire handshake_detector_stall;
  wire [7:0] handshake_generator_data;
  wire handshake_generator_issue_ack;
  wire handshake_generator_issue_nak;
  wire handshake_generator_issue_stall;
  wire handshake_generator_ready;
  wire handshake_generator_valid;
  input last;
  wire last;
  output \last$3 ;
  wire \last$3 ;
  wire low_speed_only;
  reg [2:0] microframe_number = 3'h0;
  reg [2:0] \microframe_number$next ;
  reg new_frame;
  input [7:0] payload;
  wire [7:0] payload;
  output [7:0] \payload$4 ;
  wire [7:0] \payload$4 ;
  output ready;
  wire ready;
  input \ready$5 ;
  wire \ready$5 ;
  wire [3:0] receiver_active_pid;
  wire [15:0] receiver_crc;
  wire receiver_crc_mismatch;
  wire receiver_next;
  wire receiver_packet_complete;
  wire [7:0] receiver_payload;
  wire receiver_ready_for_response;
  wire receiver_start;
  wire \receiver_start$9 ;
  wire receiver_tx_allowed;
  wire receiver_valid;
  wire reset_detected;
  wire reset_sequencer_bus_busy;
  wire reset_sequencer_bus_reset;
  wire [1:0] reset_sequencer_current_speed;
  wire [7:0] reset_sequencer_data;
  wire reset_sequencer_full_speed_only;
  wire [1:0] reset_sequencer_line_state;
  wire reset_sequencer_low_speed_only;
  wire [1:0] reset_sequencer_operating_mode;
  wire reset_sequencer_suspended;
  wire reset_sequencer_termination_select;
  wire reset_sequencer_valid;
  wire rx_activity_led;
  wire sof_detected;
  wire [1:0] speed;
  wire suspended;
  wire timer_rx_timeout;
  wire [1:0] timer_speed;
  wire timer_start;
  wire timer_tx_allowed;
  wire timer_tx_timeout;
  wire [6:0] token_detector_address;
  wire [6:0] \token_detector_address$6 ;
  wire [3:0] token_detector_endpoint;
  wire [10:0] token_detector_frame;
  wire token_detector_is_in;
  wire token_detector_is_out;
  wire token_detector_is_ping;
  wire token_detector_is_setup;
  wire token_detector_new_frame;
  wire token_detector_new_token;
  wire [3:0] token_detector_pid;
  wire token_detector_ready_for_response;
  wire [1:0] token_detector_speed;
  wire translator_busy;
  wire translator_dm_pulldown;
  wire translator_dp_pulldown;
  wire [1:0] translator_line_state;
  wire [1:0] translator_op_mode;
  wire translator_rx_active;
  wire [7:0] translator_rx_data;
  wire translator_rx_valid;
  wire translator_session_end;
  wire translator_term_select;
  wire [7:0] translator_tx_data;
  wire translator_tx_ready;
  wire translator_tx_valid;
  wire [1:0] translator_xcvr_select;
  wire [15:0] transmitter_crc;
  wire [7:0] transmitter_data;
  wire [1:0] transmitter_data_pid;
  wire transmitter_first;
  wire transmitter_last;
  wire [7:0] transmitter_payload;
  wire transmitter_ready;
  wire \transmitter_ready$8 ;
  wire transmitter_start;
  wire transmitter_valid;
  wire \transmitter_valid$7 ;
  wire tx_activity_led;
  wire [7:0] tx_multiplexer_data;
  wire tx_multiplexer_ready;
  wire tx_multiplexer_valid;
  input ulpi__clk;
  wire ulpi__clk;
  input [7:0] ulpi__data__i;
  wire [7:0] ulpi__data__i;
  output [7:0] ulpi__data__o;
  wire [7:0] ulpi__data__o;
  output ulpi__data__oe;
  wire ulpi__data__oe;
  input ulpi__dir__i;
  wire ulpi__dir__i;
  input ulpi__nxt;
  wire ulpi__nxt;
  output ulpi__rst;
  wire ulpi__rst;
  output ulpi__stp;
  wire ulpi__stp;
  output usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  input valid;
  wire valid;
  output \valid$1 ;
  wire \valid$1 ;
  wire vbus_connected;
  assign \$111  = ~  translator_session_end;
  assign \$113  = +  receiver_active_pid[3];
  assign \$115  = tx_multiplexer_valid &  translator_tx_ready;
  assign \$124  = reset_sequencer_termination_select &  connect;
  assign \$126  = token_detector_frame !=  frame_number;
  assign \$129  = microframe_number +  1'h1;
  always @(posedge usb_clk)
    address <= \address$next ;
  always @(posedge usb_clk)
    configuration <= \configuration$next ;
  always @(posedge usb_clk)
    frame_number <= \frame_number$next ;
  always @(posedge usb_clk)
    microframe_number <= \microframe_number$next ;
  USBControlEndpoint USBControlEndpoint (
    .ack(\endpoint_mux_ack$15 ),
    .\ack$1 (\endpoint_mux_ack$81 ),
    .active_config(\endpoint_mux_active_config$35 ),
    .address(\endpoint_mux_address$20 ),
    .address_changed(\endpoint_mux_address_changed$77 ),
    .config_changed(\endpoint_mux_config_changed$79 ),
    .crc(endpoint_mux_crc),
    .endpoint(\endpoint_mux_endpoint$21 ),
    .first(\endpoint_mux_first$102 ),
    .frame(\endpoint_mux_frame$24 ),
    .is_in(\endpoint_mux_is_in$26 ),
    .is_out(\endpoint_mux_is_out$27 ),
    .is_ping(\endpoint_mux_is_ping$29 ),
    .is_setup(\endpoint_mux_is_setup$28 ),
    .last(\endpoint_mux_last$105 ),
    .nak(\endpoint_mux_nak$16 ),
    .\nak$2 (\endpoint_mux_nak$85 ),
    .new_address(\endpoint_mux_new_address$78 ),
    .new_config(\endpoint_mux_new_config$80 ),
    .new_frame(\endpoint_mux_new_frame$25 ),
    .new_token(\endpoint_mux_new_token$22 ),
    .next(\endpoint_mux_next$31 ),
    .nyet(\endpoint_mux_nyet$18 ),
    .payload(\endpoint_mux_payload$32 ),
    .\payload$6 (\endpoint_mux_payload$99 ),
    .pid(\endpoint_mux_pid$19 ),
    .ready(\endpoint_mux_ready$108 ),
    .ready_for_response(\endpoint_mux_ready_for_response$23 ),
    .rx_active(translator_rx_active),
    .rx_data(translator_rx_data),
    .rx_ready_for_response(\endpoint_mux_rx_ready_for_response$33 ),
    .rx_timeout(endpoint_mux_rx_timeout),
    .rx_valid(translator_rx_valid),
    .speed(\endpoint_mux_speed$34 ),
    .stall(\endpoint_mux_stall$17 ),
    .\stall$3 (\endpoint_mux_stall$89 ),
    .start(endpoint_mux_start),
    .\start$4 (\endpoint_mux_start$92 ),
    .tx_allowed(endpoint_mux_tx_allowed),
    .tx_pid_toggle(\endpoint_mux_tx_pid_toggle$96 ),
    .tx_timeout(endpoint_mux_tx_timeout),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst),
    .valid(\endpoint_mux_valid$30 ),
    .\valid$5 (\endpoint_mux_valid$93 )
  );
  USBStreamInEndpoint USBStreamInEndpoint (
    .ack(\endpoint_mux_ack$36 ),
    .\ack$1 (\endpoint_mux_ack$82 ),
    .address(\endpoint_mux_address$41 ),
    .endpoint(\endpoint_mux_endpoint$42 ),
    .first(\endpoint_mux_first$103 ),
    .frame(\endpoint_mux_frame$45 ),
    .is_in(\endpoint_mux_is_in$47 ),
    .is_out(\endpoint_mux_is_out$48 ),
    .is_ping(\endpoint_mux_is_ping$50 ),
    .is_setup(\endpoint_mux_is_setup$49 ),
    .last(\endpoint_mux_last$106 ),
    .nak(\endpoint_mux_nak$37 ),
    .\nak$2 (\endpoint_mux_nak$86 ),
    .new_frame(\endpoint_mux_new_frame$46 ),
    .new_token(\endpoint_mux_new_token$43 ),
    .nyet(\endpoint_mux_nyet$39 ),
    .payload(\endpoint_mux_payload$100 ),
    .pid(\endpoint_mux_pid$40 ),
    .ready(\endpoint_mux_ready$109 ),
    .ready_for_response(\endpoint_mux_ready_for_response$44 ),
    .stall(\endpoint_mux_stall$38 ),
    .\stall$3 (\endpoint_mux_stall$90 ),
    .tx_pid_toggle(\endpoint_mux_tx_pid_toggle$97 ),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst),
    .valid(\endpoint_mux_valid$94 )
  );
  USBStreamInEndpoint_2831507112816 USBStreamInEndpoint_2831507112816 (
    .ack(\endpoint_mux_ack$62 ),
    .\ack$1 (\endpoint_mux_ack$84 ),
    .address(\endpoint_mux_address$67 ),
    .endpoint(\endpoint_mux_endpoint$68 ),
    .first(first),
    .\first$6 (\endpoint_mux_first$104 ),
    .frame(\endpoint_mux_frame$71 ),
    .is_in(\endpoint_mux_is_in$73 ),
    .is_out(\endpoint_mux_is_out$74 ),
    .is_ping(\endpoint_mux_is_ping$76 ),
    .is_setup(\endpoint_mux_is_setup$75 ),
    .last(last),
    .\last$7 (\endpoint_mux_last$107 ),
    .nak(\endpoint_mux_nak$63 ),
    .\nak$2 (\endpoint_mux_nak$88 ),
    .new_frame(\endpoint_mux_new_frame$72 ),
    .new_token(\endpoint_mux_new_token$69 ),
    .nyet(\endpoint_mux_nyet$65 ),
    .payload(payload),
    .\payload$5 (\endpoint_mux_payload$101 ),
    .pid(\endpoint_mux_pid$66 ),
    .ready(ready),
    .\ready$8 (\endpoint_mux_ready$110 ),
    .ready_for_response(\endpoint_mux_ready_for_response$70 ),
    .stall(\endpoint_mux_stall$64 ),
    .\stall$3 (\endpoint_mux_stall$91 ),
    .tx_pid_toggle(\endpoint_mux_tx_pid_toggle$98 ),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst),
    .valid(valid),
    .\valid$4 (\endpoint_mux_valid$95 )
  );
  USBStreamOutEndpoint USBStreamOutEndpoint (
    .ack(\endpoint_mux_ack$83 ),
    .endpoint(\endpoint_mux_endpoint$51 ),
    .first(\first$2 ),
    .is_out(\endpoint_mux_is_out$53 ),
    .is_ping(\endpoint_mux_is_ping$54 ),
    .last(\last$3 ),
    .nak(\endpoint_mux_nak$87 ),
    .next(\endpoint_mux_next$56 ),
    .payload(\payload$4 ),
    .\payload$2 (\endpoint_mux_payload$57 ),
    .ready(\ready$5 ),
    .ready_for_response(\endpoint_mux_ready_for_response$52 ),
    .rx_complete(\endpoint_mux_rx_complete$58 ),
    .rx_invalid(\endpoint_mux_rx_invalid$60 ),
    .rx_pid_toggle(\endpoint_mux_rx_pid_toggle$61 ),
    .rx_ready_for_response(\endpoint_mux_rx_ready_for_response$59 ),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst),
    .valid(\valid$1 ),
    .\valid$1 (\endpoint_mux_valid$55 )
  );
  data_crc data_crc (
    .crc(transmitter_crc),
    .\crc$2 (receiver_crc),
    .\crc$4 (data_crc_crc),
    .rx_data(data_crc_rx_data),
    .rx_valid(data_crc_rx_valid),
    .start(transmitter_start),
    .\start$1 (receiver_start),
    .\start$3 (data_crc_start),
    .tx_data(data_crc_tx_data),
    .tx_valid(data_crc_tx_valid),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst)
  );
  endpoint_mux endpoint_mux (
    .ack(endpoint_mux_ack),
    .\ack$11 (\endpoint_mux_ack$15 ),
    .\ack$3 (\endpoint_mux_ack$12 ),
    .\ack$32 (\endpoint_mux_ack$36 ),
    .\ack$58 (\endpoint_mux_ack$62 ),
    .\ack$77 (\endpoint_mux_ack$81 ),
    .\ack$78 (\endpoint_mux_ack$82 ),
    .\ack$79 (\endpoint_mux_ack$83 ),
    .\ack$80 (\endpoint_mux_ack$84 ),
    .active_address(endpoint_mux_active_address),
    .active_config(endpoint_mux_active_config),
    .\active_config$31 (\endpoint_mux_active_config$35 ),
    .address(endpoint_mux_address),
    .\address$16 (\endpoint_mux_address$20 ),
    .\address$37 (\endpoint_mux_address$41 ),
    .\address$63 (\endpoint_mux_address$67 ),
    .address_changed(endpoint_mux_address_changed),
    .\address_changed$73 (\endpoint_mux_address_changed$77 ),
    .config_changed(endpoint_mux_config_changed),
    .\config_changed$75 (\endpoint_mux_config_changed$79 ),
    .crc(data_crc_crc),
    .\crc$7 (endpoint_mux_crc),
    .endpoint(endpoint_mux_endpoint),
    .\endpoint$17 (\endpoint_mux_endpoint$21 ),
    .\endpoint$38 (\endpoint_mux_endpoint$42 ),
    .\endpoint$47 (\endpoint_mux_endpoint$51 ),
    .\endpoint$64 (\endpoint_mux_endpoint$68 ),
    .first(endpoint_mux_first),
    .\first$100 (\endpoint_mux_first$103 ),
    .\first$101 (\endpoint_mux_first$104 ),
    .\first$99 (\endpoint_mux_first$102 ),
    .frame(endpoint_mux_frame),
    .\frame$20 (\endpoint_mux_frame$24 ),
    .\frame$41 (\endpoint_mux_frame$45 ),
    .\frame$67 (\endpoint_mux_frame$71 ),
    .is_in(endpoint_mux_is_in),
    .\is_in$22 (\endpoint_mux_is_in$26 ),
    .\is_in$43 (\endpoint_mux_is_in$47 ),
    .\is_in$69 (\endpoint_mux_is_in$73 ),
    .is_out(endpoint_mux_is_out),
    .\is_out$23 (\endpoint_mux_is_out$27 ),
    .\is_out$44 (\endpoint_mux_is_out$48 ),
    .\is_out$49 (\endpoint_mux_is_out$53 ),
    .\is_out$70 (\endpoint_mux_is_out$74 ),
    .is_ping(endpoint_mux_is_ping),
    .\is_ping$25 (\endpoint_mux_is_ping$29 ),
    .\is_ping$46 (\endpoint_mux_is_ping$50 ),
    .\is_ping$50 (\endpoint_mux_is_ping$54 ),
    .\is_ping$72 (\endpoint_mux_is_ping$76 ),
    .is_setup(endpoint_mux_is_setup),
    .\is_setup$24 (\endpoint_mux_is_setup$28 ),
    .\is_setup$45 (\endpoint_mux_is_setup$49 ),
    .\is_setup$71 (\endpoint_mux_is_setup$75 ),
    .last(endpoint_mux_last),
    .\last$102 (\endpoint_mux_last$105 ),
    .\last$103 (\endpoint_mux_last$106 ),
    .\last$104 (\endpoint_mux_last$107 ),
    .nak(endpoint_mux_nak),
    .\nak$12 (\endpoint_mux_nak$16 ),
    .\nak$33 (\endpoint_mux_nak$37 ),
    .\nak$4 (\endpoint_mux_nak$13 ),
    .\nak$59 (\endpoint_mux_nak$63 ),
    .\nak$81 (\endpoint_mux_nak$85 ),
    .\nak$82 (\endpoint_mux_nak$86 ),
    .\nak$83 (\endpoint_mux_nak$87 ),
    .\nak$84 (\endpoint_mux_nak$88 ),
    .new_address(endpoint_mux_new_address),
    .\new_address$74 (\endpoint_mux_new_address$78 ),
    .new_config(endpoint_mux_new_config),
    .\new_config$76 (\endpoint_mux_new_config$80 ),
    .new_frame(endpoint_mux_new_frame),
    .\new_frame$21 (\endpoint_mux_new_frame$25 ),
    .\new_frame$42 (\endpoint_mux_new_frame$46 ),
    .\new_frame$68 (\endpoint_mux_new_frame$72 ),
    .new_token(endpoint_mux_new_token),
    .\new_token$18 (\endpoint_mux_new_token$22 ),
    .\new_token$39 (\endpoint_mux_new_token$43 ),
    .\new_token$65 (\endpoint_mux_new_token$69 ),
    .next(endpoint_mux_next),
    .\next$27 (\endpoint_mux_next$31 ),
    .\next$52 (\endpoint_mux_next$56 ),
    .nyet(endpoint_mux_nyet),
    .\nyet$14 (\endpoint_mux_nyet$18 ),
    .\nyet$35 (\endpoint_mux_nyet$39 ),
    .\nyet$61 (\endpoint_mux_nyet$65 ),
    .payload(endpoint_mux_payload),
    .\payload$2 (\endpoint_mux_payload$11 ),
    .\payload$28 (\endpoint_mux_payload$32 ),
    .\payload$53 (\endpoint_mux_payload$57 ),
    .\payload$96 (\endpoint_mux_payload$99 ),
    .\payload$97 (\endpoint_mux_payload$100 ),
    .\payload$98 (\endpoint_mux_payload$101 ),
    .pid(endpoint_mux_pid),
    .\pid$15 (\endpoint_mux_pid$19 ),
    .\pid$36 (\endpoint_mux_pid$40 ),
    .\pid$62 (\endpoint_mux_pid$66 ),
    .ready(endpoint_mux_ready),
    .\ready$105 (\endpoint_mux_ready$108 ),
    .\ready$106 (\endpoint_mux_ready$109 ),
    .\ready$107 (\endpoint_mux_ready$110 ),
    .ready_for_response(endpoint_mux_ready_for_response),
    .\ready_for_response$19 (\endpoint_mux_ready_for_response$23 ),
    .\ready_for_response$40 (\endpoint_mux_ready_for_response$44 ),
    .\ready_for_response$48 (\endpoint_mux_ready_for_response$52 ),
    .\ready_for_response$66 (\endpoint_mux_ready_for_response$70 ),
    .rx_complete(endpoint_mux_rx_complete),
    .\rx_complete$54 (\endpoint_mux_rx_complete$58 ),
    .rx_invalid(endpoint_mux_rx_invalid),
    .\rx_invalid$56 (\endpoint_mux_rx_invalid$60 ),
    .rx_pid_toggle(endpoint_mux_rx_pid_toggle),
    .\rx_pid_toggle$57 (\endpoint_mux_rx_pid_toggle$61 ),
    .rx_ready_for_response(endpoint_mux_rx_ready_for_response),
    .\rx_ready_for_response$29 (\endpoint_mux_rx_ready_for_response$33 ),
    .\rx_ready_for_response$55 (\endpoint_mux_rx_ready_for_response$59 ),
    .rx_timeout(timer_rx_timeout),
    .\rx_timeout$10 (endpoint_mux_rx_timeout),
    .speed(endpoint_mux_speed),
    .\speed$30 (\endpoint_mux_speed$34 ),
    .stall(endpoint_mux_stall),
    .\stall$13 (\endpoint_mux_stall$17 ),
    .\stall$34 (\endpoint_mux_stall$38 ),
    .\stall$5 (\endpoint_mux_stall$14 ),
    .\stall$60 (\endpoint_mux_stall$64 ),
    .\stall$85 (\endpoint_mux_stall$89 ),
    .\stall$86 (\endpoint_mux_stall$90 ),
    .\stall$87 (\endpoint_mux_stall$91 ),
    .start(data_crc_start),
    .\start$6 (timer_start),
    .\start$88 (endpoint_mux_start),
    .\start$89 (\endpoint_mux_start$92 ),
    .tx_allowed(timer_tx_allowed),
    .\tx_allowed$8 (endpoint_mux_tx_allowed),
    .tx_pid_toggle(endpoint_mux_tx_pid_toggle),
    .\tx_pid_toggle$93 (\endpoint_mux_tx_pid_toggle$96 ),
    .\tx_pid_toggle$94 (\endpoint_mux_tx_pid_toggle$97 ),
    .\tx_pid_toggle$95 (\endpoint_mux_tx_pid_toggle$98 ),
    .tx_timeout(timer_tx_timeout),
    .\tx_timeout$9 (endpoint_mux_tx_timeout),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst),
    .valid(endpoint_mux_valid),
    .\valid$1 (\endpoint_mux_valid$10 ),
    .\valid$26 (\endpoint_mux_valid$30 ),
    .\valid$51 (\endpoint_mux_valid$55 ),
    .\valid$90 (\endpoint_mux_valid$93 ),
    .\valid$91 (\endpoint_mux_valid$94 ),
    .\valid$92 (\endpoint_mux_valid$95 )
  );
  handshake_detector handshake_detector (
    .ack(handshake_detector_ack),
    .nak(handshake_detector_nak),
    .nyet(handshake_detector_nyet),
    .rx_active(translator_rx_active),
    .rx_data(translator_rx_data),
    .rx_valid(translator_rx_valid),
    .stall(handshake_detector_stall),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst)
  );
  handshake_generator handshake_generator (
    .data(handshake_generator_data),
    .issue_ack(handshake_generator_issue_ack),
    .issue_nak(handshake_generator_issue_nak),
    .issue_stall(handshake_generator_issue_stall),
    .ready(handshake_generator_ready),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst),
    .valid(handshake_generator_valid)
  );
  receiver receiver (
    .active_pid(receiver_active_pid),
    .crc(receiver_crc),
    .crc_mismatch(receiver_crc_mismatch),
    .next(receiver_next),
    .packet_complete(receiver_packet_complete),
    .payload(receiver_payload),
    .ready_for_response(receiver_ready_for_response),
    .rx_active(translator_rx_active),
    .rx_data(translator_rx_data),
    .rx_valid(translator_rx_valid),
    .start(receiver_start),
    .\start$1 (\receiver_start$9 ),
    .tx_allowed(receiver_tx_allowed),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst),
    .valid(receiver_valid)
  );
  reset_sequencer reset_sequencer (
    .bus_busy(reset_sequencer_bus_busy),
    .bus_reset(reset_sequencer_bus_reset),
    .current_speed(reset_sequencer_current_speed),
    .data(reset_sequencer_data),
    .full_speed_only(1'h0),
    .line_state(reset_sequencer_line_state),
    .low_speed_only(1'h0),
    .operating_mode(reset_sequencer_operating_mode),
    .suspended(reset_sequencer_suspended),
    .termination_select(reset_sequencer_termination_select),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst),
    .valid(reset_sequencer_valid)
  );
  \timer$1  timer (
    .rx_timeout(timer_rx_timeout),
    .speed(timer_speed),
    .start(\receiver_start$9 ),
    .\start$1 (timer_start),
    .tx_allowed(receiver_tx_allowed),
    .\tx_allowed$2 (timer_tx_allowed),
    .tx_timeout(timer_tx_timeout),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst)
  );
  token_detector token_detector (
    .address(token_detector_address),
    .\address$1 (\token_detector_address$6 ),
    .endpoint(token_detector_endpoint),
    .frame(token_detector_frame),
    .is_in(token_detector_is_in),
    .is_out(token_detector_is_out),
    .is_ping(token_detector_is_ping),
    .is_setup(token_detector_is_setup),
    .new_frame(token_detector_new_frame),
    .new_token(token_detector_new_token),
    .pid(token_detector_pid),
    .ready_for_response(token_detector_ready_for_response),
    .rx_active(translator_rx_active),
    .rx_data(translator_rx_data),
    .rx_valid(translator_rx_valid),
    .speed(token_detector_speed),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst)
  );
  translator translator (
    .busy(translator_busy),
    .dm_pulldown(1'h0),
    .dp_pulldown(1'h0),
    .line_state(translator_line_state),
    .op_mode(translator_op_mode),
    .rx_active(translator_rx_active),
    .rx_data(translator_rx_data),
    .rx_valid(translator_rx_valid),
    .session_end(translator_session_end),
    .term_select(translator_term_select),
    .tx_data(translator_tx_data),
    .tx_ready(translator_tx_ready),
    .tx_valid(translator_tx_valid),
    .ulpi__clk(ulpi__clk),
    .ulpi__data__i(ulpi__data__i),
    .ulpi__data__o(ulpi__data__o),
    .ulpi__data__oe(ulpi__data__oe),
    .ulpi__dir__i(ulpi__dir__i),
    .ulpi__nxt(ulpi__nxt),
    .ulpi__rst(ulpi__rst),
    .ulpi__stp(ulpi__stp),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst),
    .xcvr_select(translator_xcvr_select)
  );
  transmitter transmitter (
    .crc(transmitter_crc),
    .data(transmitter_data),
    .data_pid(transmitter_data_pid),
    .first(transmitter_first),
    .last(transmitter_last),
    .payload(transmitter_payload),
    .ready(transmitter_ready),
    .\ready$2 (\transmitter_ready$8 ),
    .start(transmitter_start),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst),
    .valid(transmitter_valid),
    .\valid$1 (\transmitter_valid$7 )
  );
  tx_multiplexer tx_multiplexer (
    .data(tx_multiplexer_data),
    .\data$2 (reset_sequencer_data),
    .\data$3 (transmitter_data),
    .\data$7 (handshake_generator_data),
    .ready(tx_multiplexer_ready),
    .\ready$5 (\transmitter_ready$8 ),
    .\ready$8 (handshake_generator_ready),
    .valid(tx_multiplexer_valid),
    .\valid$1 (reset_sequencer_valid),
    .\valid$4 (\transmitter_valid$7 ),
    .\valid$6 (handshake_generator_valid)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$36 ) begin end
    \address$next  = address;
    casez (endpoint_mux_address_changed)
      1'h1:
          \address$next  = endpoint_mux_new_address;
    endcase
    casez (reset_sequencer_bus_reset)
      1'h1:
          \address$next  = 7'h00;
    endcase
    casez (usb_rst)
      1'h1:
          \address$next  = 7'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$36 ) begin end
    \configuration$next  = configuration;
    casez (endpoint_mux_config_changed)
      1'h1:
          \configuration$next  = endpoint_mux_new_config;
    endcase
    casez (reset_sequencer_bus_reset)
      1'h1:
          \configuration$next  = 8'h00;
    endcase
    casez (usb_rst)
      1'h1:
          \configuration$next  = 8'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$36 ) begin end
    \frame_number$next  = frame_number;
    casez (token_detector_new_frame)
      1'h1:
          \frame_number$next  = token_detector_frame;
    endcase
    casez (usb_rst)
      1'h1:
          \frame_number$next  = 11'h000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$36 ) begin end
    new_frame = 1'h0;
    casez (token_detector_new_frame)
      1'h1:
          new_frame = \$126 ;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$36 ) begin end
    \microframe_number$next  = microframe_number;
    casez (token_detector_new_frame)
      1'h1:
          casez (new_frame)
            1'h1:
                \microframe_number$next  = 3'h0;
            default:
                \microframe_number$next  = \$129 [2:0];
          endcase
    endcase
    casez (usb_rst)
      1'h1:
          \microframe_number$next  = 3'h0;
    endcase
  end
  assign \$117  = \$120 ;
  assign \$128  = \$129 ;
  assign low_speed_only = 1'h0;
  assign full_speed_only = 1'h0;
  assign rx_activity_led = translator_rx_valid;
  assign tx_activity_led = tx_multiplexer_valid;
  assign reset_detected = reset_sequencer_bus_reset;
  assign sof_detected = token_detector_new_frame;
  assign suspended = reset_sequencer_suspended;
  assign speed = reset_sequencer_current_speed;
  assign translator_term_select = \$124 ;
  assign translator_xcvr_select = reset_sequencer_current_speed;
  assign translator_op_mode = reset_sequencer_operating_mode;
  assign reset_sequencer_full_speed_only = \$122 ;
  assign reset_sequencer_low_speed_only = \$120 [0];
  assign translator_dp_pulldown = 1'h0;
  assign translator_dm_pulldown = 1'h0;
  assign data_crc_tx_data = tx_multiplexer_data;
  assign data_crc_tx_valid = \$115 ;
  assign tx_multiplexer_ready = translator_tx_ready;
  assign translator_tx_valid = tx_multiplexer_valid;
  assign translator_tx_data = tx_multiplexer_data;
  assign transmitter_data_pid = endpoint_mux_tx_pid_toggle;
  assign handshake_generator_issue_stall = \endpoint_mux_stall$14 ;
  assign handshake_generator_issue_nak = \endpoint_mux_nak$13 ;
  assign handshake_generator_issue_ack = \endpoint_mux_ack$12 ;
  assign endpoint_mux_ready = transmitter_ready;
  assign transmitter_payload = \endpoint_mux_payload$11 ;
  assign transmitter_last = endpoint_mux_last;
  assign transmitter_first = endpoint_mux_first;
  assign transmitter_valid = \endpoint_mux_valid$10 ;
  assign endpoint_mux_rx_pid_toggle = \$113 ;
  assign endpoint_mux_rx_ready_for_response = receiver_ready_for_response;
  assign endpoint_mux_rx_invalid = receiver_crc_mismatch;
  assign endpoint_mux_rx_complete = receiver_packet_complete;
  assign endpoint_mux_payload = receiver_payload;
  assign endpoint_mux_next = receiver_next;
  assign endpoint_mux_valid = receiver_valid;
  assign endpoint_mux_active_address = address;
  assign endpoint_mux_active_config = configuration;
  assign endpoint_mux_speed = speed;
  assign endpoint_mux_nyet = handshake_detector_nyet;
  assign endpoint_mux_stall = handshake_detector_stall;
  assign endpoint_mux_nak = handshake_detector_nak;
  assign endpoint_mux_ack = handshake_detector_ack;
  assign endpoint_mux_is_ping = token_detector_is_ping;
  assign endpoint_mux_is_setup = token_detector_is_setup;
  assign endpoint_mux_is_out = token_detector_is_out;
  assign endpoint_mux_is_in = token_detector_is_in;
  assign endpoint_mux_new_frame = token_detector_new_frame;
  assign endpoint_mux_frame = token_detector_frame;
  assign endpoint_mux_ready_for_response = token_detector_ready_for_response;
  assign endpoint_mux_new_token = token_detector_new_token;
  assign endpoint_mux_endpoint = token_detector_endpoint;
  assign endpoint_mux_address = \token_detector_address$6 ;
  assign endpoint_mux_pid = token_detector_pid;
  assign timer_speed = speed;
  assign token_detector_speed = speed;
  assign data_crc_rx_valid = translator_rx_valid;
  assign data_crc_rx_data = translator_rx_data;
  assign token_detector_address = address;
  assign reset_sequencer_line_state = translator_line_state;
  assign vbus_connected = \$111 ;
  assign reset_sequencer_bus_busy = translator_busy;
  assign \$118  = 2'h0;
  assign \$120  = 2'h0;
  assign \$122  = 1'h0;
endmodule
module usb_serial(ulpi__data__o, ulpi__data__oe, ulpi__clk, ulpi__nxt, ulpi__stp, ulpi__dir__i, ulpi__rst, tx__valid, tx__ready, tx__first, tx__last, tx__payload, rx__valid, rx__ready, rx__first, rx__last, rx__payload, usb_clk, usb_rst, ulpi__data__i);
  output rx__first;
  wire rx__first;
  output rx__last;
  wire rx__last;
  output [7:0] rx__payload;
  wire [7:0] rx__payload;
  input rx__ready;
  wire rx__ready;
  output rx__valid;
  wire rx__valid;
  input tx__first;
  wire tx__first;
  input tx__last;
  wire tx__last;
  input [7:0] tx__payload;
  wire [7:0] tx__payload;
  output tx__ready;
  wire tx__ready;
  input tx__valid;
  wire tx__valid;
  input ulpi__clk;
  wire ulpi__clk;
  input [7:0] ulpi__data__i;
  wire [7:0] ulpi__data__i;
  output [7:0] ulpi__data__o;
  wire [7:0] ulpi__data__o;
  output ulpi__data__oe;
  wire ulpi__data__oe;
  input ulpi__dir__i;
  wire ulpi__dir__i;
  input ulpi__nxt;
  wire ulpi__nxt;
  output ulpi__rst;
  wire ulpi__rst;
  output ulpi__stp;
  wire ulpi__stp;
  output usb_clk;
  wire usb_clk;
  input usb_rst;
  wire usb_rst;
  wire usb_serial_device_connect;
  wire usb_serial_device_first;
  wire \usb_serial_device_first$2 ;
  wire usb_serial_device_last;
  wire \usb_serial_device_last$3 ;
  wire [7:0] usb_serial_device_payload;
  wire [7:0] \usb_serial_device_payload$4 ;
  wire usb_serial_device_ready;
  wire \usb_serial_device_ready$5 ;
  wire usb_serial_device_valid;
  wire \usb_serial_device_valid$1 ;
  usb_serial_device usb_serial_device (
    .connect(1'h1),
    .first(usb_serial_device_first),
    .\first$2 (\usb_serial_device_first$2 ),
    .last(usb_serial_device_last),
    .\last$3 (\usb_serial_device_last$3 ),
    .payload(usb_serial_device_payload),
    .\payload$4 (\usb_serial_device_payload$4 ),
    .ready(usb_serial_device_ready),
    .\ready$5 (\usb_serial_device_ready$5 ),
    .ulpi__clk(ulpi__clk),
    .ulpi__data__i(ulpi__data__i),
    .ulpi__data__o(ulpi__data__o),
    .ulpi__data__oe(ulpi__data__oe),
    .ulpi__dir__i(ulpi__dir__i),
    .ulpi__nxt(ulpi__nxt),
    .ulpi__rst(ulpi__rst),
    .ulpi__stp(ulpi__stp),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst),
    .valid(usb_serial_device_valid),
    .\valid$1 (\usb_serial_device_valid$1 )
  );
  assign \usb_serial_device_ready$5  = rx__ready;
  assign rx__payload = \usb_serial_device_payload$4 ;
  assign rx__last = \usb_serial_device_last$3 ;
  assign rx__first = \usb_serial_device_first$2 ;
  assign rx__valid = \usb_serial_device_valid$1 ;
  assign tx__ready = usb_serial_device_ready;
  assign usb_serial_device_payload = tx__payload;
  assign usb_serial_device_last = tx__last;
  assign usb_serial_device_first = tx__first;
  assign usb_serial_device_valid = tx__valid;
  assign usb_serial_device_connect = 1'h1;
endmodule
module usb_serial_device(valid, first, last, payload, ready, \valid$1 , \first$2 , \last$3 , \payload$4 , \ready$5 , usb_rst, usb_clk, ulpi__clk, ulpi__rst, ulpi__data__oe, ulpi__dir__i, ulpi__nxt, ulpi__data__i, ulpi__data__o, ulpi__stp, connect
);
  input connect;
  wire connect;
  input first;
  wire first;
  output \first$2 ;
  wire \first$2 ;
  input last;
  wire last;
  output \last$3 ;
  wire \last$3 ;
  input [7:0] payload;
  wire [7:0] payload;
  output [7:0] \payload$4 ;
  wire [7:0] \payload$4 ;
  output ready;
  wire ready;
  input \ready$5 ;
  wire \ready$5 ;
  input ulpi__clk;
  wire ulpi__clk;
  input [7:0] ulpi__data__i;
  wire [7:0] ulpi__data__i;
  output [7:0] ulpi__data__o;
  wire [7:0] ulpi__data__o;
  output ulpi__data__oe;
  wire ulpi__data__oe;
  input ulpi__dir__i;
  wire ulpi__dir__i;
  input ulpi__nxt;
  wire ulpi__nxt;
  output ulpi__rst;
  wire ulpi__rst;
  output ulpi__stp;
  wire ulpi__stp;
  output usb_clk;
  wire usb_clk;
  wire usb_connect;
  wire usb_first;
  wire \usb_first$7 ;
  wire usb_last;
  wire \usb_last$8 ;
  wire [7:0] usb_payload;
  wire [7:0] \usb_payload$9 ;
  wire usb_ready;
  wire \usb_ready$10 ;
  input usb_rst;
  wire usb_rst;
  wire usb_valid;
  wire \usb_valid$6 ;
  input valid;
  wire valid;
  output \valid$1 ;
  wire \valid$1 ;
  usb usb (
    .connect(usb_connect),
    .first(usb_first),
    .\first$2 (\usb_first$7 ),
    .last(usb_last),
    .\last$3 (\usb_last$8 ),
    .payload(usb_payload),
    .\payload$4 (\usb_payload$9 ),
    .ready(usb_ready),
    .\ready$5 (\usb_ready$10 ),
    .ulpi__clk(ulpi__clk),
    .ulpi__data__i(ulpi__data__i),
    .ulpi__data__o(ulpi__data__o),
    .ulpi__data__oe(ulpi__data__oe),
    .ulpi__dir__i(ulpi__dir__i),
    .ulpi__nxt(ulpi__nxt),
    .ulpi__rst(ulpi__rst),
    .ulpi__stp(ulpi__stp),
    .usb_clk(usb_clk),
    .usb_rst(usb_rst),
    .valid(usb_valid),
    .\valid$1 (\usb_valid$6 )
  );
  assign usb_connect = connect;
  assign \usb_ready$10  = \ready$5 ;
  assign \payload$4  = \usb_payload$9 ;
  assign \last$3  = \usb_last$8 ;
  assign \first$2  = \usb_first$7 ;
  assign \valid$1  = \usb_valid$6 ;
  assign ready = usb_ready;
  assign usb_payload = payload;
  assign usb_last = last;
  assign usb_first = first;
  assign usb_valid = valid;
endmodule
