module ddr3_top (
	input fifo_clk,    // Clock
	input video_clk,

	
	
);

endmodule